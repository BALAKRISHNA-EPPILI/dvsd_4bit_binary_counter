* NGSPICE file created from dvsd_4bit_binary_counter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt dvsd_4bit_binary_counter VGND VPWR clk out[0] out[1] out[2] out[3] reset updown
X_49_ _49_/CLK _49_/D VGND VGND VPWR VPWR _49_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_48_ _49_/CLK _48_/D VGND VGND VPWR VPWR _48_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/CLK _47_/D VGND VGND VPWR VPWR _47_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ _47_/CLK _46_/D VGND VGND VPWR VPWR _46_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_29_ _46_/Q _47_/Q VGND VGND VPWR VPWR _35_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28_ _46_/Q _47_/Q VGND VGND VPWR VPWR _32_/B sky130_fd_sc_hd__or2_1
X_45_ _38_/X _40_/X _45_/S VGND VGND VPWR VPWR _45_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_44_ _33_/X _36_/X _45_/S VGND VGND VPWR VPWR _44_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/A VGND VGND VPWR VPWR _27_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_43_ _31_/A _31_/Y _45_/S VGND VGND VPWR VPWR _43_/X sky130_fd_sc_hd__mux2_1
X_26_ _46_/Q VGND VGND VPWR VPWR _27_/A sky130_fd_sc_hd__inv_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_42_ _27_/A _27_/X _45_/S VGND VGND VPWR VPWR _42_/X sky130_fd_sc_hd__mux2_1
X_25_ _41_/A _42_/X VGND VGND VPWR VPWR _46_/D sky130_fd_sc_hd__nor2b_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24_ _41_/A _43_/X VGND VGND VPWR VPWR _47_/D sky130_fd_sc_hd__nor2b_1
X_41_ _41_/A _45_/X VGND VGND VPWR VPWR _49_/D sky130_fd_sc_hd__nor2b_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_40_ _48_/Q _35_/Y _37_/Y _39_/X VGND VGND VPWR VPWR _40_/X sky130_fd_sc_hd__a31o_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23_ _41_/A _44_/X VGND VGND VPWR VPWR _48_/D sky130_fd_sc_hd__nor2b_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 reset VGND VGND VPWR VPWR _41_/A sky130_fd_sc_hd__buf_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 updown VGND VGND VPWR VPWR _45_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _49_/CLK sky130_fd_sc_hd__clkbuf_16
X_39_ _34_/Y _35_/A _49_/Q VGND VGND VPWR VPWR _39_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ _37_/Y _32_/X _37_/Y _32_/X VGND VGND VPWR VPWR _38_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_37_ _49_/Q VGND VGND VPWR VPWR _37_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36_ _34_/Y _35_/A _48_/Q _35_/Y VGND VGND VPWR VPWR _36_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35_ _35_/A VGND VGND VPWR VPWR _35_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34_ _48_/Q VGND VGND VPWR VPWR _34_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33_ _48_/Q _32_/B _32_/X VGND VGND VPWR VPWR _33_/X sky130_fd_sc_hd__a21bo_1
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _47_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ _48_/Q _32_/B VGND VGND VPWR VPWR _32_/X sky130_fd_sc_hd__or2_1
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ _31_/A VGND VGND VPWR VPWR _31_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30_ _32_/B _35_/A VGND VGND VPWR VPWR _31_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput3 _46_/Q VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput4 _47_/Q VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput5 _48_/Q VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput6 _49_/Q VGND VGND VPWR VPWR out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

