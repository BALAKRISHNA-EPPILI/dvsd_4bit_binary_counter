magic
tech sky130A
magscale 1 2
timestamp 1629458243
<< viali >>
rect 2881 11781 2915 11815
rect 3065 11713 3099 11747
rect 9505 11713 9539 11747
rect 9321 11509 9355 11543
rect 3985 10013 4019 10047
rect 6561 10013 6595 10047
rect 3801 9945 3835 9979
rect 4169 9945 4203 9979
rect 6377 9945 6411 9979
rect 6745 9945 6779 9979
rect 3056 9605 3090 9639
rect 8493 9605 8527 9639
rect 1961 9537 1995 9571
rect 4905 9537 4939 9571
rect 2789 9469 2823 9503
rect 4813 9469 4847 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 1869 9333 1903 9367
rect 4169 9333 4203 9367
rect 4629 9333 4663 9367
rect 7021 9333 7055 9367
rect 5549 9129 5583 9163
rect 3157 8993 3191 9027
rect 4261 8993 4295 9027
rect 6929 8993 6963 9027
rect 3249 8925 3283 8959
rect 4353 8925 4387 8959
rect 4724 8925 4758 8959
rect 6662 8925 6696 8959
rect 7573 8925 7607 8959
rect 7389 8857 7423 8891
rect 7757 8857 7791 8891
rect 4721 8789 4755 8823
rect 4905 8789 4939 8823
rect 4261 8585 4295 8619
rect 4629 8585 4663 8619
rect 4721 8517 4755 8551
rect 5457 8517 5491 8551
rect 7766 8517 7800 8551
rect 2421 8449 2455 8483
rect 2688 8449 2722 8483
rect 5641 8449 5675 8483
rect 4905 8381 4939 8415
rect 8033 8381 8067 8415
rect 3801 8313 3835 8347
rect 5825 8245 5859 8279
rect 6653 8245 6687 8279
rect 2881 8041 2915 8075
rect 6285 8041 6319 8075
rect 7481 8041 7515 8075
rect 4629 7905 4663 7939
rect 5365 7905 5399 7939
rect 6929 7905 6963 7939
rect 8125 7905 8159 7939
rect 3065 7837 3099 7871
rect 5457 7837 5491 7871
rect 3249 7769 3283 7803
rect 4353 7769 4387 7803
rect 5181 7769 5215 7803
rect 5825 7769 5859 7803
rect 7849 7769 7883 7803
rect 3985 7701 4019 7735
rect 4445 7701 4479 7735
rect 6653 7701 6687 7735
rect 6745 7701 6779 7735
rect 7941 7701 7975 7735
rect 3065 7497 3099 7531
rect 4813 7497 4847 7531
rect 7297 7497 7331 7531
rect 9137 7497 9171 7531
rect 4353 7429 4387 7463
rect 7849 7429 7883 7463
rect 4997 7361 5031 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 7205 7361 7239 7395
rect 5273 7157 5307 7191
rect 6469 7157 6503 7191
rect 4905 6953 4939 6987
rect 6377 6953 6411 6987
rect 8953 6953 8987 6987
rect 4997 6817 5031 6851
rect 5457 6817 5491 6851
rect 7021 6817 7055 6851
rect 3985 6749 4019 6783
rect 4721 6749 4755 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 6929 6749 6963 6783
rect 9137 6749 9171 6783
rect 4537 6681 4571 6715
rect 3893 6613 3927 6647
rect 4997 6409 5031 6443
rect 4905 6273 4939 6307
rect 10333 2533 10367 2567
rect 1961 2397 1995 2431
rect 6929 2397 6963 2431
rect 1777 2329 1811 2363
rect 6745 2329 6779 2363
rect 10517 2329 10551 2363
<< metal1 >>
rect 1104 11994 11316 12016
rect 1104 11942 4386 11994
rect 4438 11942 4450 11994
rect 4502 11942 4514 11994
rect 4566 11942 4578 11994
rect 4630 11942 7790 11994
rect 7842 11942 7854 11994
rect 7906 11942 7918 11994
rect 7970 11942 7982 11994
rect 8034 11942 11316 11994
rect 1104 11920 11316 11942
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 2869 11815 2927 11821
rect 2869 11812 2881 11815
rect 2832 11784 2881 11812
rect 2832 11772 2838 11784
rect 2869 11781 2881 11784
rect 2915 11781 2927 11815
rect 2869 11775 2927 11781
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9272 11716 9505 11744
rect 9272 11704 9278 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9306 11540 9312 11552
rect 9267 11512 9312 11540
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 1104 11450 11316 11472
rect 1104 11398 2684 11450
rect 2736 11398 2748 11450
rect 2800 11398 2812 11450
rect 2864 11398 2876 11450
rect 2928 11398 6088 11450
rect 6140 11398 6152 11450
rect 6204 11398 6216 11450
rect 6268 11398 6280 11450
rect 6332 11398 9492 11450
rect 9544 11398 9556 11450
rect 9608 11398 9620 11450
rect 9672 11398 9684 11450
rect 9736 11398 11316 11450
rect 1104 11376 11316 11398
rect 1104 10906 11316 10928
rect 1104 10854 4386 10906
rect 4438 10854 4450 10906
rect 4502 10854 4514 10906
rect 4566 10854 4578 10906
rect 4630 10854 7790 10906
rect 7842 10854 7854 10906
rect 7906 10854 7918 10906
rect 7970 10854 7982 10906
rect 8034 10854 11316 10906
rect 1104 10832 11316 10854
rect 1104 10362 11316 10384
rect 1104 10310 2684 10362
rect 2736 10310 2748 10362
rect 2800 10310 2812 10362
rect 2864 10310 2876 10362
rect 2928 10310 6088 10362
rect 6140 10310 6152 10362
rect 6204 10310 6216 10362
rect 6268 10310 6280 10362
rect 6332 10310 9492 10362
rect 9544 10310 9556 10362
rect 9608 10310 9620 10362
rect 9672 10310 9684 10362
rect 9736 10310 11316 10362
rect 1104 10288 11316 10310
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 3384 10016 3985 10044
rect 3384 10004 3390 10016
rect 3973 10013 3985 10016
rect 4019 10044 4031 10047
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 4019 10016 6561 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 6549 10013 6561 10016
rect 6595 10044 6607 10047
rect 7558 10044 7564 10056
rect 6595 10016 7564 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7558 10004 7564 10016
rect 7616 10044 7622 10056
rect 9306 10044 9312 10056
rect 7616 10016 9312 10044
rect 7616 10004 7622 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 3786 9976 3792 9988
rect 3747 9948 3792 9976
rect 3786 9936 3792 9948
rect 3844 9936 3850 9988
rect 4154 9976 4160 9988
rect 4115 9948 4160 9976
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 6365 9979 6423 9985
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 6454 9976 6460 9988
rect 6411 9948 6460 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6696 9948 6745 9976
rect 6696 9936 6702 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 1104 9818 11316 9840
rect 1104 9766 4386 9818
rect 4438 9766 4450 9818
rect 4502 9766 4514 9818
rect 4566 9766 4578 9818
rect 4630 9766 7790 9818
rect 7842 9766 7854 9818
rect 7906 9766 7918 9818
rect 7970 9766 7982 9818
rect 8034 9766 11316 9818
rect 1104 9744 11316 9766
rect 3044 9639 3102 9645
rect 3044 9605 3056 9639
rect 3090 9636 3102 9639
rect 3786 9636 3792 9648
rect 3090 9608 3792 9636
rect 3090 9605 3102 9608
rect 3044 9599 3102 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 8478 9636 8484 9648
rect 8439 9608 8484 9636
rect 8478 9596 8484 9608
rect 8536 9596 8542 9648
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 4893 9571 4951 9577
rect 1995 9540 4660 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2792 9364 2820 9463
rect 4632 9432 4660 9540
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5166 9568 5172 9580
rect 4939 9540 5172 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 4798 9500 4804 9512
rect 4759 9472 4804 9500
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4982 9500 4988 9512
rect 4943 9472 4988 9500
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5132 9472 5177 9500
rect 5132 9460 5138 9472
rect 5534 9432 5540 9444
rect 4632 9404 5540 9432
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 3142 9364 3148 9376
rect 2792 9336 3148 9364
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4246 9364 4252 9376
rect 4203 9336 4252 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4706 9364 4712 9376
rect 4663 9336 4712 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6972 9336 7021 9364
rect 6972 9324 6978 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 1104 9274 11316 9296
rect 1104 9222 2684 9274
rect 2736 9222 2748 9274
rect 2800 9222 2812 9274
rect 2864 9222 2876 9274
rect 2928 9222 6088 9274
rect 6140 9222 6152 9274
rect 6204 9222 6216 9274
rect 6268 9222 6280 9274
rect 6332 9222 9492 9274
rect 9544 9222 9556 9274
rect 9608 9222 9620 9274
rect 9672 9222 9684 9274
rect 9736 9222 11316 9274
rect 1104 9200 11316 9222
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 3191 8996 4261 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 4249 8993 4261 8996
rect 4295 9024 4307 9027
rect 6917 9027 6975 9033
rect 4295 8996 4476 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3108 8928 3249 8956
rect 3108 8916 3114 8928
rect 3237 8925 3249 8928
rect 3283 8956 3295 8959
rect 4341 8959 4399 8965
rect 3283 8928 4292 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 4264 8900 4292 8928
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4448 8956 4476 8996
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 8386 9024 8392 9036
rect 6963 8996 8392 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 4712 8959 4770 8965
rect 4712 8956 4724 8959
rect 4448 8928 4724 8956
rect 4341 8919 4399 8925
rect 4712 8925 4724 8928
rect 4758 8956 4770 8959
rect 4798 8956 4804 8968
rect 4758 8928 4804 8956
rect 4758 8925 4770 8928
rect 4712 8919 4770 8925
rect 4246 8848 4252 8900
rect 4304 8848 4310 8900
rect 4356 8820 4384 8919
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 6638 8916 6644 8968
rect 6696 8965 6702 8968
rect 6696 8956 6708 8965
rect 7558 8956 7564 8968
rect 6696 8928 6741 8956
rect 7519 8928 7564 8956
rect 6696 8919 6708 8928
rect 6696 8916 6702 8919
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 5350 8888 5356 8900
rect 4724 8860 5356 8888
rect 4724 8829 4752 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 7374 8888 7380 8900
rect 7335 8860 7380 8888
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 7650 8848 7656 8900
rect 7708 8888 7714 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7708 8860 7757 8888
rect 7708 8848 7714 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 4709 8823 4767 8829
rect 4709 8820 4721 8823
rect 4356 8792 4721 8820
rect 4709 8789 4721 8792
rect 4755 8789 4767 8823
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4709 8783 4767 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 1104 8730 11316 8752
rect 1104 8678 4386 8730
rect 4438 8678 4450 8730
rect 4502 8678 4514 8730
rect 4566 8678 4578 8730
rect 4630 8678 7790 8730
rect 7842 8678 7854 8730
rect 7906 8678 7918 8730
rect 7970 8678 7982 8730
rect 8034 8678 11316 8730
rect 1104 8656 11316 8678
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4212 8588 4261 8616
rect 4212 8576 4218 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4890 8616 4896 8628
rect 4663 8588 4896 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 3142 8548 3148 8560
rect 2424 8520 3148 8548
rect 2424 8489 2452 8520
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 4706 8548 4712 8560
rect 4667 8520 4712 8548
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 5445 8551 5503 8557
rect 5445 8517 5457 8551
rect 5491 8548 5503 8551
rect 5534 8548 5540 8560
rect 5491 8520 5540 8548
rect 5491 8517 5503 8520
rect 5445 8511 5503 8517
rect 5534 8508 5540 8520
rect 5592 8548 5598 8560
rect 6546 8548 6552 8560
rect 5592 8520 6552 8548
rect 5592 8508 5598 8520
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 7754 8551 7812 8557
rect 7754 8548 7766 8551
rect 7708 8520 7766 8548
rect 7708 8508 7714 8520
rect 7754 8517 7766 8520
rect 7800 8517 7812 8551
rect 7754 8511 7812 8517
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2676 8483 2734 8489
rect 2676 8449 2688 8483
rect 2722 8480 2734 8483
rect 3050 8480 3056 8492
rect 2722 8452 3056 8480
rect 2722 8449 2734 8452
rect 2676 8443 2734 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 5675 8452 6684 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 4890 8412 4896 8424
rect 4851 8384 4896 8412
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8344 3847 8347
rect 4982 8344 4988 8356
rect 3835 8316 4988 8344
rect 3835 8313 3847 8316
rect 3789 8307 3847 8313
rect 4982 8304 4988 8316
rect 5040 8304 5046 8356
rect 5810 8276 5816 8288
rect 5771 8248 5816 8276
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 6656 8285 6684 8452
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8386 8412 8392 8424
rect 8067 8384 8392 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 6730 8276 6736 8288
rect 6687 8248 6736 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 1104 8186 11316 8208
rect 1104 8134 2684 8186
rect 2736 8134 2748 8186
rect 2800 8134 2812 8186
rect 2864 8134 2876 8186
rect 2928 8134 6088 8186
rect 6140 8134 6152 8186
rect 6204 8134 6216 8186
rect 6268 8134 6280 8186
rect 6332 8134 9492 8186
rect 9544 8134 9556 8186
rect 9608 8134 9620 8186
rect 9672 8134 9684 8186
rect 9736 8134 11316 8186
rect 1104 8112 11316 8134
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3050 8072 3056 8084
rect 2915 8044 3056 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 6273 8075 6331 8081
rect 6273 8041 6285 8075
rect 6319 8072 6331 8075
rect 6454 8072 6460 8084
rect 6319 8044 6460 8072
rect 6319 8041 6331 8044
rect 6273 8035 6331 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7432 8044 7481 8072
rect 7432 8032 7438 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 4890 8004 4896 8016
rect 4632 7976 4896 8004
rect 4632 7945 4660 7976
rect 4890 7964 4896 7976
rect 4948 8004 4954 8016
rect 4948 7976 6960 8004
rect 4948 7964 4954 7976
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5810 7936 5816 7948
rect 5399 7908 5816 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6932 7945 6960 7976
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 6963 7908 8125 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 8113 7905 8125 7908
rect 8159 7936 8171 7939
rect 10318 7936 10324 7948
rect 8159 7908 10324 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3326 7868 3332 7880
rect 3099 7840 3332 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5040 7840 5457 7868
rect 5040 7828 5046 7840
rect 5445 7837 5457 7840
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7769 3295 7803
rect 3237 7763 3295 7769
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 5169 7803 5227 7809
rect 5169 7800 5181 7803
rect 4387 7772 5181 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 5169 7769 5181 7772
rect 5215 7769 5227 7803
rect 5169 7763 5227 7769
rect 3252 7732 3280 7763
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 5408 7772 5825 7800
rect 5408 7760 5414 7772
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 5813 7763 5871 7769
rect 7837 7803 7895 7809
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 8294 7800 8300 7812
rect 7883 7772 8300 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 8294 7760 8300 7772
rect 8352 7800 8358 7812
rect 9122 7800 9128 7812
rect 8352 7772 9128 7800
rect 8352 7760 8358 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3252 7704 3985 7732
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4798 7732 4804 7744
rect 4479 7704 4804 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6733 7735 6791 7741
rect 6733 7701 6745 7735
rect 6779 7732 6791 7735
rect 7006 7732 7012 7744
rect 6779 7704 7012 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8938 7732 8944 7744
rect 7975 7704 8944 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 1104 7642 11316 7664
rect 1104 7590 4386 7642
rect 4438 7590 4450 7642
rect 4502 7590 4514 7642
rect 4566 7590 4578 7642
rect 4630 7590 7790 7642
rect 7842 7590 7854 7642
rect 7906 7590 7918 7642
rect 7970 7590 7982 7642
rect 8034 7590 11316 7642
rect 1104 7568 11316 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3142 7528 3148 7540
rect 3099 7500 3148 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4798 7528 4804 7540
rect 4759 7500 4804 7528
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 8294 7528 8300 7540
rect 7331 7500 8300 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8444 7500 9137 7528
rect 8444 7488 8450 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 6914 7460 6920 7472
rect 4387 7432 6920 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 6914 7420 6920 7432
rect 6972 7460 6978 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 6972 7432 7849 7460
rect 6972 7420 6978 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 4982 7392 4988 7404
rect 4856 7364 4988 7392
rect 4856 7352 4862 7364
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5166 7392 5172 7404
rect 5123 7364 5172 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5350 7392 5356 7404
rect 5311 7364 5356 7392
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6365 7355 6423 7361
rect 6380 7324 6408 7355
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 7190 7392 7196 7404
rect 7151 7364 7196 7392
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 6730 7324 6736 7336
rect 6380 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7324 6794 7336
rect 7208 7324 7236 7352
rect 6788 7296 7236 7324
rect 6788 7284 6794 7296
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4948 7160 5273 7188
rect 4948 7148 4954 7160
rect 5261 7157 5273 7160
rect 5307 7188 5319 7191
rect 6454 7188 6460 7200
rect 5307 7160 6460 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 1104 7098 11316 7120
rect 1104 7046 2684 7098
rect 2736 7046 2748 7098
rect 2800 7046 2812 7098
rect 2864 7046 2876 7098
rect 2928 7046 6088 7098
rect 6140 7046 6152 7098
rect 6204 7046 6216 7098
rect 6268 7046 6280 7098
rect 6332 7046 9492 7098
rect 9544 7046 9556 7098
rect 9608 7046 9620 7098
rect 9672 7046 9684 7098
rect 9736 7046 11316 7098
rect 1104 7024 11316 7046
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 6638 6984 6644 6996
rect 6411 6956 6644 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 8938 6984 8944 6996
rect 8899 6956 8944 6984
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 4908 6916 4936 6944
rect 4816 6888 4936 6916
rect 4816 6848 4844 6888
rect 4982 6848 4988 6860
rect 3988 6820 4844 6848
rect 4895 6820 4988 6848
rect 3988 6789 4016 6820
rect 4982 6808 4988 6820
rect 5040 6848 5046 6860
rect 5350 6848 5356 6860
rect 5040 6820 5356 6848
rect 5040 6808 5046 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 7006 6848 7012 6860
rect 5500 6820 5545 6848
rect 6967 6820 7012 6848
rect 5500 6808 5506 6820
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4304 6752 4721 6780
rect 4304 6740 4310 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5629 6783 5687 6789
rect 5629 6780 5641 6783
rect 4948 6752 5641 6780
rect 4948 6740 4954 6752
rect 5629 6749 5641 6752
rect 5675 6749 5687 6783
rect 5810 6780 5816 6792
rect 5771 6752 5816 6780
rect 5629 6743 5687 6749
rect 5810 6740 5816 6752
rect 5868 6780 5874 6792
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5868 6752 6285 6780
rect 5868 6740 5874 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6273 6743 6331 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6696 6752 6929 6780
rect 6696 6740 6702 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 6917 6743 6975 6749
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 4525 6715 4583 6721
rect 4525 6681 4537 6715
rect 4571 6712 4583 6715
rect 5074 6712 5080 6724
rect 4571 6684 5080 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 5074 6672 5080 6684
rect 5132 6672 5138 6724
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 5166 6644 5172 6656
rect 3927 6616 5172 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 1104 6554 11316 6576
rect 1104 6502 4386 6554
rect 4438 6502 4450 6554
rect 4502 6502 4514 6554
rect 4566 6502 4578 6554
rect 4630 6502 7790 6554
rect 7842 6502 7854 6554
rect 7906 6502 7918 6554
rect 7970 6502 7982 6554
rect 8034 6502 11316 6554
rect 1104 6480 11316 6502
rect 4982 6440 4988 6452
rect 4943 6412 4988 6440
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 1104 6010 11316 6032
rect 1104 5958 2684 6010
rect 2736 5958 2748 6010
rect 2800 5958 2812 6010
rect 2864 5958 2876 6010
rect 2928 5958 6088 6010
rect 6140 5958 6152 6010
rect 6204 5958 6216 6010
rect 6268 5958 6280 6010
rect 6332 5958 9492 6010
rect 9544 5958 9556 6010
rect 9608 5958 9620 6010
rect 9672 5958 9684 6010
rect 9736 5958 11316 6010
rect 1104 5936 11316 5958
rect 1104 5466 11316 5488
rect 1104 5414 4386 5466
rect 4438 5414 4450 5466
rect 4502 5414 4514 5466
rect 4566 5414 4578 5466
rect 4630 5414 7790 5466
rect 7842 5414 7854 5466
rect 7906 5414 7918 5466
rect 7970 5414 7982 5466
rect 8034 5414 11316 5466
rect 1104 5392 11316 5414
rect 1104 4922 11316 4944
rect 1104 4870 2684 4922
rect 2736 4870 2748 4922
rect 2800 4870 2812 4922
rect 2864 4870 2876 4922
rect 2928 4870 6088 4922
rect 6140 4870 6152 4922
rect 6204 4870 6216 4922
rect 6268 4870 6280 4922
rect 6332 4870 9492 4922
rect 9544 4870 9556 4922
rect 9608 4870 9620 4922
rect 9672 4870 9684 4922
rect 9736 4870 11316 4922
rect 1104 4848 11316 4870
rect 1104 4378 11316 4400
rect 1104 4326 4386 4378
rect 4438 4326 4450 4378
rect 4502 4326 4514 4378
rect 4566 4326 4578 4378
rect 4630 4326 7790 4378
rect 7842 4326 7854 4378
rect 7906 4326 7918 4378
rect 7970 4326 7982 4378
rect 8034 4326 11316 4378
rect 1104 4304 11316 4326
rect 1104 3834 11316 3856
rect 1104 3782 2684 3834
rect 2736 3782 2748 3834
rect 2800 3782 2812 3834
rect 2864 3782 2876 3834
rect 2928 3782 6088 3834
rect 6140 3782 6152 3834
rect 6204 3782 6216 3834
rect 6268 3782 6280 3834
rect 6332 3782 9492 3834
rect 9544 3782 9556 3834
rect 9608 3782 9620 3834
rect 9672 3782 9684 3834
rect 9736 3782 11316 3834
rect 1104 3760 11316 3782
rect 1104 3290 11316 3312
rect 1104 3238 4386 3290
rect 4438 3238 4450 3290
rect 4502 3238 4514 3290
rect 4566 3238 4578 3290
rect 4630 3238 7790 3290
rect 7842 3238 7854 3290
rect 7906 3238 7918 3290
rect 7970 3238 7982 3290
rect 8034 3238 11316 3290
rect 1104 3216 11316 3238
rect 1104 2746 11316 2768
rect 1104 2694 2684 2746
rect 2736 2694 2748 2746
rect 2800 2694 2812 2746
rect 2864 2694 2876 2746
rect 2928 2694 6088 2746
rect 6140 2694 6152 2746
rect 6204 2694 6216 2746
rect 6268 2694 6280 2746
rect 6332 2694 9492 2746
rect 9544 2694 9556 2746
rect 9608 2694 9620 2746
rect 9672 2694 9684 2746
rect 9736 2694 11316 2746
rect 1104 2672 11316 2694
rect 10318 2564 10324 2576
rect 10279 2536 10324 2564
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 4890 2428 4896 2440
rect 1995 2400 4896 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7190 2428 7196 2440
rect 6963 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 72 2332 1777 2360
rect 72 2320 78 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 6270 2320 6276 2372
rect 6328 2360 6334 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6328 2332 6745 2360
rect 6328 2320 6334 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 10502 2360 10508 2372
rect 10463 2332 10508 2360
rect 6733 2323 6791 2329
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 1104 2202 11316 2224
rect 1104 2150 4386 2202
rect 4438 2150 4450 2202
rect 4502 2150 4514 2202
rect 4566 2150 4578 2202
rect 4630 2150 7790 2202
rect 7842 2150 7854 2202
rect 7906 2150 7918 2202
rect 7970 2150 7982 2202
rect 8034 2150 11316 2202
rect 1104 2128 11316 2150
<< via1 >>
rect 4386 11942 4438 11994
rect 4450 11942 4502 11994
rect 4514 11942 4566 11994
rect 4578 11942 4630 11994
rect 7790 11942 7842 11994
rect 7854 11942 7906 11994
rect 7918 11942 7970 11994
rect 7982 11942 8034 11994
rect 2780 11772 2832 11824
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 9220 11704 9272 11756
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 2684 11398 2736 11450
rect 2748 11398 2800 11450
rect 2812 11398 2864 11450
rect 2876 11398 2928 11450
rect 6088 11398 6140 11450
rect 6152 11398 6204 11450
rect 6216 11398 6268 11450
rect 6280 11398 6332 11450
rect 9492 11398 9544 11450
rect 9556 11398 9608 11450
rect 9620 11398 9672 11450
rect 9684 11398 9736 11450
rect 4386 10854 4438 10906
rect 4450 10854 4502 10906
rect 4514 10854 4566 10906
rect 4578 10854 4630 10906
rect 7790 10854 7842 10906
rect 7854 10854 7906 10906
rect 7918 10854 7970 10906
rect 7982 10854 8034 10906
rect 2684 10310 2736 10362
rect 2748 10310 2800 10362
rect 2812 10310 2864 10362
rect 2876 10310 2928 10362
rect 6088 10310 6140 10362
rect 6152 10310 6204 10362
rect 6216 10310 6268 10362
rect 6280 10310 6332 10362
rect 9492 10310 9544 10362
rect 9556 10310 9608 10362
rect 9620 10310 9672 10362
rect 9684 10310 9736 10362
rect 3332 10004 3384 10056
rect 7564 10004 7616 10056
rect 9312 10004 9364 10056
rect 3792 9979 3844 9988
rect 3792 9945 3801 9979
rect 3801 9945 3835 9979
rect 3835 9945 3844 9979
rect 3792 9936 3844 9945
rect 4160 9979 4212 9988
rect 4160 9945 4169 9979
rect 4169 9945 4203 9979
rect 4203 9945 4212 9979
rect 4160 9936 4212 9945
rect 6460 9936 6512 9988
rect 6644 9936 6696 9988
rect 4386 9766 4438 9818
rect 4450 9766 4502 9818
rect 4514 9766 4566 9818
rect 4578 9766 4630 9818
rect 7790 9766 7842 9818
rect 7854 9766 7906 9818
rect 7918 9766 7970 9818
rect 7982 9766 8034 9818
rect 3792 9596 3844 9648
rect 8484 9639 8536 9648
rect 8484 9605 8493 9639
rect 8493 9605 8527 9639
rect 8527 9605 8536 9639
rect 8484 9596 8536 9605
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 5172 9528 5224 9580
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5540 9392 5592 9444
rect 3148 9324 3200 9376
rect 4252 9324 4304 9376
rect 4712 9324 4764 9376
rect 6920 9324 6972 9376
rect 2684 9222 2736 9274
rect 2748 9222 2800 9274
rect 2812 9222 2864 9274
rect 2876 9222 2928 9274
rect 6088 9222 6140 9274
rect 6152 9222 6204 9274
rect 6216 9222 6268 9274
rect 6280 9222 6332 9274
rect 9492 9222 9544 9274
rect 9556 9222 9608 9274
rect 9620 9222 9672 9274
rect 9684 9222 9736 9274
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 3056 8916 3108 8968
rect 8392 8984 8444 9036
rect 4252 8848 4304 8900
rect 4804 8916 4856 8968
rect 6644 8959 6696 8968
rect 6644 8925 6662 8959
rect 6662 8925 6696 8959
rect 7564 8959 7616 8968
rect 6644 8916 6696 8925
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 5356 8848 5408 8900
rect 7380 8891 7432 8900
rect 7380 8857 7389 8891
rect 7389 8857 7423 8891
rect 7423 8857 7432 8891
rect 7380 8848 7432 8857
rect 7656 8848 7708 8900
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 4386 8678 4438 8730
rect 4450 8678 4502 8730
rect 4514 8678 4566 8730
rect 4578 8678 4630 8730
rect 7790 8678 7842 8730
rect 7854 8678 7906 8730
rect 7918 8678 7970 8730
rect 7982 8678 8034 8730
rect 4160 8576 4212 8628
rect 4896 8576 4948 8628
rect 3148 8508 3200 8560
rect 4712 8551 4764 8560
rect 4712 8517 4721 8551
rect 4721 8517 4755 8551
rect 4755 8517 4764 8551
rect 4712 8508 4764 8517
rect 5540 8508 5592 8560
rect 6552 8508 6604 8560
rect 7656 8508 7708 8560
rect 3056 8440 3108 8492
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 4988 8304 5040 8356
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 8392 8372 8444 8424
rect 6736 8236 6788 8288
rect 2684 8134 2736 8186
rect 2748 8134 2800 8186
rect 2812 8134 2864 8186
rect 2876 8134 2928 8186
rect 6088 8134 6140 8186
rect 6152 8134 6204 8186
rect 6216 8134 6268 8186
rect 6280 8134 6332 8186
rect 9492 8134 9544 8186
rect 9556 8134 9608 8186
rect 9620 8134 9672 8186
rect 9684 8134 9736 8186
rect 3056 8032 3108 8084
rect 6460 8032 6512 8084
rect 7380 8032 7432 8084
rect 4896 7964 4948 8016
rect 5816 7896 5868 7948
rect 10324 7896 10376 7948
rect 3332 7828 3384 7880
rect 4988 7828 5040 7880
rect 5356 7760 5408 7812
rect 8300 7760 8352 7812
rect 9128 7760 9180 7812
rect 4804 7692 4856 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7012 7692 7064 7744
rect 8944 7692 8996 7744
rect 4386 7590 4438 7642
rect 4450 7590 4502 7642
rect 4514 7590 4566 7642
rect 4578 7590 4630 7642
rect 7790 7590 7842 7642
rect 7854 7590 7906 7642
rect 7918 7590 7970 7642
rect 7982 7590 8034 7642
rect 3148 7488 3200 7540
rect 4804 7531 4856 7540
rect 4804 7497 4813 7531
rect 4813 7497 4847 7531
rect 4847 7497 4856 7531
rect 4804 7488 4856 7497
rect 8300 7488 8352 7540
rect 8392 7488 8444 7540
rect 6920 7420 6972 7472
rect 4804 7352 4856 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5172 7352 5224 7404
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 6736 7284 6788 7336
rect 4896 7148 4948 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 2684 7046 2736 7098
rect 2748 7046 2800 7098
rect 2812 7046 2864 7098
rect 2876 7046 2928 7098
rect 6088 7046 6140 7098
rect 6152 7046 6204 7098
rect 6216 7046 6268 7098
rect 6280 7046 6332 7098
rect 9492 7046 9544 7098
rect 9556 7046 9608 7098
rect 9620 7046 9672 7098
rect 9684 7046 9736 7098
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 6644 6944 6696 6996
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5356 6808 5408 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 7012 6851 7064 6860
rect 5448 6808 5500 6817
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 4252 6740 4304 6792
rect 4896 6740 4948 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6644 6740 6696 6792
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 5080 6672 5132 6724
rect 5172 6604 5224 6656
rect 4386 6502 4438 6554
rect 4450 6502 4502 6554
rect 4514 6502 4566 6554
rect 4578 6502 4630 6554
rect 7790 6502 7842 6554
rect 7854 6502 7906 6554
rect 7918 6502 7970 6554
rect 7982 6502 8034 6554
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 2684 5958 2736 6010
rect 2748 5958 2800 6010
rect 2812 5958 2864 6010
rect 2876 5958 2928 6010
rect 6088 5958 6140 6010
rect 6152 5958 6204 6010
rect 6216 5958 6268 6010
rect 6280 5958 6332 6010
rect 9492 5958 9544 6010
rect 9556 5958 9608 6010
rect 9620 5958 9672 6010
rect 9684 5958 9736 6010
rect 4386 5414 4438 5466
rect 4450 5414 4502 5466
rect 4514 5414 4566 5466
rect 4578 5414 4630 5466
rect 7790 5414 7842 5466
rect 7854 5414 7906 5466
rect 7918 5414 7970 5466
rect 7982 5414 8034 5466
rect 2684 4870 2736 4922
rect 2748 4870 2800 4922
rect 2812 4870 2864 4922
rect 2876 4870 2928 4922
rect 6088 4870 6140 4922
rect 6152 4870 6204 4922
rect 6216 4870 6268 4922
rect 6280 4870 6332 4922
rect 9492 4870 9544 4922
rect 9556 4870 9608 4922
rect 9620 4870 9672 4922
rect 9684 4870 9736 4922
rect 4386 4326 4438 4378
rect 4450 4326 4502 4378
rect 4514 4326 4566 4378
rect 4578 4326 4630 4378
rect 7790 4326 7842 4378
rect 7854 4326 7906 4378
rect 7918 4326 7970 4378
rect 7982 4326 8034 4378
rect 2684 3782 2736 3834
rect 2748 3782 2800 3834
rect 2812 3782 2864 3834
rect 2876 3782 2928 3834
rect 6088 3782 6140 3834
rect 6152 3782 6204 3834
rect 6216 3782 6268 3834
rect 6280 3782 6332 3834
rect 9492 3782 9544 3834
rect 9556 3782 9608 3834
rect 9620 3782 9672 3834
rect 9684 3782 9736 3834
rect 4386 3238 4438 3290
rect 4450 3238 4502 3290
rect 4514 3238 4566 3290
rect 4578 3238 4630 3290
rect 7790 3238 7842 3290
rect 7854 3238 7906 3290
rect 7918 3238 7970 3290
rect 7982 3238 8034 3290
rect 2684 2694 2736 2746
rect 2748 2694 2800 2746
rect 2812 2694 2864 2746
rect 2876 2694 2928 2746
rect 6088 2694 6140 2746
rect 6152 2694 6204 2746
rect 6216 2694 6268 2746
rect 6280 2694 6332 2746
rect 9492 2694 9544 2746
rect 9556 2694 9608 2746
rect 9620 2694 9672 2746
rect 9684 2694 9736 2746
rect 10324 2567 10376 2576
rect 10324 2533 10333 2567
rect 10333 2533 10367 2567
rect 10367 2533 10376 2567
rect 10324 2524 10376 2533
rect 4896 2388 4948 2440
rect 7196 2388 7248 2440
rect 20 2320 72 2372
rect 6276 2320 6328 2372
rect 10508 2363 10560 2372
rect 10508 2329 10517 2363
rect 10517 2329 10551 2363
rect 10551 2329 10560 2363
rect 10508 2320 10560 2329
rect 4386 2150 4438 2202
rect 4450 2150 4502 2202
rect 4514 2150 4566 2202
rect 4578 2150 4630 2202
rect 7790 2150 7842 2202
rect 7854 2150 7906 2202
rect 7918 2150 7970 2202
rect 7982 2150 8034 2202
<< metal2 >>
rect 2778 13779 2834 14579
rect 9218 13779 9274 14579
rect 2792 11830 2820 13779
rect 4360 11996 4656 12016
rect 4416 11994 4440 11996
rect 4496 11994 4520 11996
rect 4576 11994 4600 11996
rect 4438 11942 4440 11994
rect 4502 11942 4514 11994
rect 4576 11942 4578 11994
rect 4416 11940 4440 11942
rect 4496 11940 4520 11942
rect 4576 11940 4600 11942
rect 4360 11920 4656 11940
rect 7764 11996 8060 12016
rect 7820 11994 7844 11996
rect 7900 11994 7924 11996
rect 7980 11994 8004 11996
rect 7842 11942 7844 11994
rect 7906 11942 7918 11994
rect 7980 11942 7982 11994
rect 7820 11940 7844 11942
rect 7900 11940 7924 11942
rect 7980 11940 8004 11942
rect 7764 11920 8060 11940
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 9232 11762 9260 13779
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 2658 11452 2954 11472
rect 2714 11450 2738 11452
rect 2794 11450 2818 11452
rect 2874 11450 2898 11452
rect 2736 11398 2738 11450
rect 2800 11398 2812 11450
rect 2874 11398 2876 11450
rect 2714 11396 2738 11398
rect 2794 11396 2818 11398
rect 2874 11396 2898 11398
rect 2658 11376 2954 11396
rect 2658 10364 2954 10384
rect 2714 10362 2738 10364
rect 2794 10362 2818 10364
rect 2874 10362 2898 10364
rect 2736 10310 2738 10362
rect 2800 10310 2812 10362
rect 2874 10310 2876 10362
rect 2714 10308 2738 10310
rect 2794 10308 2818 10310
rect 2874 10308 2898 10310
rect 2658 10288 2954 10308
rect 1860 9376 1912 9382
rect 1858 9344 1860 9353
rect 1912 9344 1914 9353
rect 1858 9279 1914 9288
rect 2658 9276 2954 9296
rect 2714 9274 2738 9276
rect 2794 9274 2818 9276
rect 2874 9274 2898 9276
rect 2736 9222 2738 9274
rect 2800 9222 2812 9274
rect 2874 9222 2876 9274
rect 2714 9220 2738 9222
rect 2794 9220 2818 9222
rect 2874 9220 2898 9222
rect 2658 9200 2954 9220
rect 3068 8974 3096 11698
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 6062 11452 6358 11472
rect 6118 11450 6142 11452
rect 6198 11450 6222 11452
rect 6278 11450 6302 11452
rect 6140 11398 6142 11450
rect 6204 11398 6216 11450
rect 6278 11398 6280 11450
rect 6118 11396 6142 11398
rect 6198 11396 6222 11398
rect 6278 11396 6302 11398
rect 6062 11376 6358 11396
rect 4360 10908 4656 10928
rect 4416 10906 4440 10908
rect 4496 10906 4520 10908
rect 4576 10906 4600 10908
rect 4438 10854 4440 10906
rect 4502 10854 4514 10906
rect 4576 10854 4578 10906
rect 4416 10852 4440 10854
rect 4496 10852 4520 10854
rect 4576 10852 4600 10854
rect 4360 10832 4656 10852
rect 7764 10908 8060 10928
rect 7820 10906 7844 10908
rect 7900 10906 7924 10908
rect 7980 10906 8004 10908
rect 7842 10854 7844 10906
rect 7906 10854 7918 10906
rect 7980 10854 7982 10906
rect 7820 10852 7844 10854
rect 7900 10852 7924 10854
rect 7980 10852 8004 10854
rect 7764 10832 8060 10852
rect 6062 10364 6358 10384
rect 6118 10362 6142 10364
rect 6198 10362 6222 10364
rect 6278 10362 6302 10364
rect 6140 10310 6142 10362
rect 6204 10310 6216 10362
rect 6278 10310 6280 10362
rect 6118 10308 6142 10310
rect 6198 10308 6222 10310
rect 6278 10308 6302 10310
rect 6062 10288 6358 10308
rect 9324 10062 9352 11494
rect 9466 11452 9762 11472
rect 9522 11450 9546 11452
rect 9602 11450 9626 11452
rect 9682 11450 9706 11452
rect 9544 11398 9546 11450
rect 9608 11398 9620 11450
rect 9682 11398 9684 11450
rect 9522 11396 9546 11398
rect 9602 11396 9626 11398
rect 9682 11396 9706 11398
rect 9466 11376 9762 11396
rect 9466 10364 9762 10384
rect 9522 10362 9546 10364
rect 9602 10362 9626 10364
rect 9682 10362 9706 10364
rect 9544 10310 9546 10362
rect 9608 10310 9620 10362
rect 9682 10310 9684 10362
rect 9522 10308 9546 10310
rect 9602 10308 9626 10310
rect 9682 10308 9706 10310
rect 9466 10288 9762 10308
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3160 8566 3188 9318
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2658 8188 2954 8208
rect 2714 8186 2738 8188
rect 2794 8186 2818 8188
rect 2874 8186 2898 8188
rect 2736 8134 2738 8186
rect 2800 8134 2812 8186
rect 2874 8134 2876 8186
rect 2714 8132 2738 8134
rect 2794 8132 2818 8134
rect 2874 8132 2898 8134
rect 2658 8112 2954 8132
rect 3068 8090 3096 8434
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3160 7546 3188 8502
rect 3344 7886 3372 9998
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 3804 9654 3832 9930
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 4172 8634 4200 9930
rect 4360 9820 4656 9840
rect 4416 9818 4440 9820
rect 4496 9818 4520 9820
rect 4576 9818 4600 9820
rect 4438 9766 4440 9818
rect 4502 9766 4514 9818
rect 4576 9766 4578 9818
rect 4416 9764 4440 9766
rect 4496 9764 4520 9766
rect 4576 9764 4600 9766
rect 4360 9744 4656 9764
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4264 8906 4292 9318
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2658 7100 2954 7120
rect 2714 7098 2738 7100
rect 2794 7098 2818 7100
rect 2874 7098 2898 7100
rect 2736 7046 2738 7098
rect 2800 7046 2812 7098
rect 2874 7046 2876 7098
rect 2714 7044 2738 7046
rect 2794 7044 2818 7046
rect 2874 7044 2898 7046
rect 2658 7024 2954 7044
rect 4264 6798 4292 8842
rect 4360 8732 4656 8752
rect 4416 8730 4440 8732
rect 4496 8730 4520 8732
rect 4576 8730 4600 8732
rect 4438 8678 4440 8730
rect 4502 8678 4514 8730
rect 4576 8678 4578 8730
rect 4416 8676 4440 8678
rect 4496 8676 4520 8678
rect 4576 8676 4600 8678
rect 4360 8656 4656 8676
rect 4724 8566 4752 9318
rect 4816 8974 4844 9454
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8634 4936 8774
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 8022 4936 8366
rect 5000 8362 5028 9454
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 5000 7886 5028 8298
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4360 7644 4656 7664
rect 4416 7642 4440 7644
rect 4496 7642 4520 7644
rect 4576 7642 4600 7644
rect 4438 7590 4440 7642
rect 4502 7590 4514 7642
rect 4576 7590 4578 7642
rect 4416 7588 4440 7590
rect 4496 7588 4520 7590
rect 4576 7588 4600 7590
rect 4360 7568 4656 7588
rect 4816 7546 4844 7686
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5000 7410 5028 7822
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4816 6882 4844 7346
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 7002 4936 7142
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4816 6854 4936 6882
rect 4908 6798 4936 6854
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4360 6556 4656 6576
rect 4416 6554 4440 6556
rect 4496 6554 4520 6556
rect 4576 6554 4600 6556
rect 4438 6502 4440 6554
rect 4502 6502 4514 6554
rect 4576 6502 4578 6554
rect 4416 6500 4440 6502
rect 4496 6500 4520 6502
rect 4576 6500 4600 6502
rect 4360 6480 4656 6500
rect 4908 6322 4936 6734
rect 5000 6458 5028 6802
rect 5092 6730 5120 9454
rect 5184 7410 5212 9522
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 9178 5580 9386
rect 6062 9276 6358 9296
rect 6118 9274 6142 9276
rect 6198 9274 6222 9276
rect 6278 9274 6302 9276
rect 6140 9222 6142 9274
rect 6204 9222 6216 9274
rect 6278 9222 6280 9274
rect 6118 9220 6142 9222
rect 6198 9220 6222 9222
rect 6278 9220 6302 9222
rect 6062 9200 6358 9220
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 7818 5396 8842
rect 5552 8566 5580 9114
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7954 5856 8230
rect 6062 8188 6358 8208
rect 6118 8186 6142 8188
rect 6198 8186 6222 8188
rect 6278 8186 6302 8188
rect 6140 8134 6142 8186
rect 6204 8134 6216 8186
rect 6278 8134 6280 8186
rect 6118 8132 6142 8134
rect 6198 8132 6222 8134
rect 6278 8132 6302 8134
rect 6062 8112 6358 8132
rect 6472 8090 6500 9930
rect 6656 8974 6684 9930
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5368 7698 5396 7754
rect 5368 7670 5488 7698
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5184 6662 5212 7346
rect 5368 6866 5396 7346
rect 5460 6866 5488 7670
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5828 6798 5856 7890
rect 6564 7410 6592 8502
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6062 7100 6358 7120
rect 6118 7098 6142 7100
rect 6198 7098 6222 7100
rect 6278 7098 6302 7100
rect 6140 7046 6142 7098
rect 6204 7046 6216 7098
rect 6278 7046 6280 7098
rect 6118 7044 6142 7046
rect 6198 7044 6222 7046
rect 6278 7044 6302 7046
rect 6062 7024 6358 7044
rect 6472 6798 6500 7142
rect 6656 7002 6684 7686
rect 6748 7342 6776 8230
rect 6932 7478 6960 9318
rect 7576 8974 7604 9998
rect 8482 9888 8538 9897
rect 7764 9820 8060 9840
rect 8482 9823 8538 9832
rect 7820 9818 7844 9820
rect 7900 9818 7924 9820
rect 7980 9818 8004 9820
rect 7842 9766 7844 9818
rect 7906 9766 7918 9818
rect 7980 9766 7982 9818
rect 7820 9764 7844 9766
rect 7900 9764 7924 9766
rect 7980 9764 8004 9766
rect 7764 9744 8060 9764
rect 8496 9654 8524 9823
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 9466 9276 9762 9296
rect 9522 9274 9546 9276
rect 9602 9274 9626 9276
rect 9682 9274 9706 9276
rect 9544 9222 9546 9274
rect 9608 9222 9620 9274
rect 9682 9222 9684 9274
rect 9522 9220 9546 9222
rect 9602 9220 9626 9222
rect 9682 9220 9706 9222
rect 9466 9200 9762 9220
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7392 8090 7420 8842
rect 7668 8566 7696 8842
rect 7764 8732 8060 8752
rect 7820 8730 7844 8732
rect 7900 8730 7924 8732
rect 7980 8730 8004 8732
rect 7842 8678 7844 8730
rect 7906 8678 7918 8730
rect 7980 8678 7982 8730
rect 7820 8676 7844 8678
rect 7900 8676 7924 8678
rect 7980 8676 8004 8678
rect 7764 8656 8060 8676
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 8404 8430 8432 8978
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6656 6798 6684 6938
rect 7024 6866 7052 7686
rect 7764 7644 8060 7664
rect 7820 7642 7844 7644
rect 7900 7642 7924 7644
rect 7980 7642 8004 7644
rect 7842 7590 7844 7642
rect 7906 7590 7918 7642
rect 7980 7590 7982 7642
rect 7820 7588 7844 7590
rect 7900 7588 7924 7590
rect 7980 7588 8004 7590
rect 7764 7568 8060 7588
rect 8312 7546 8340 7754
rect 8404 7546 8432 8366
rect 9466 8188 9762 8208
rect 9522 8186 9546 8188
rect 9602 8186 9626 8188
rect 9682 8186 9706 8188
rect 9544 8134 9546 8186
rect 9608 8134 9620 8186
rect 9682 8134 9684 8186
rect 9522 8132 9546 8134
rect 9602 8132 9626 8134
rect 9682 8132 9706 8134
rect 9466 8112 9762 8132
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 2658 6012 2954 6032
rect 2714 6010 2738 6012
rect 2794 6010 2818 6012
rect 2874 6010 2898 6012
rect 2736 5958 2738 6010
rect 2800 5958 2812 6010
rect 2874 5958 2876 6010
rect 2714 5956 2738 5958
rect 2794 5956 2818 5958
rect 2874 5956 2898 5958
rect 2658 5936 2954 5956
rect 4360 5468 4656 5488
rect 4416 5466 4440 5468
rect 4496 5466 4520 5468
rect 4576 5466 4600 5468
rect 4438 5414 4440 5466
rect 4502 5414 4514 5466
rect 4576 5414 4578 5466
rect 4416 5412 4440 5414
rect 4496 5412 4520 5414
rect 4576 5412 4600 5414
rect 4360 5392 4656 5412
rect 2658 4924 2954 4944
rect 2714 4922 2738 4924
rect 2794 4922 2818 4924
rect 2874 4922 2898 4924
rect 2736 4870 2738 4922
rect 2800 4870 2812 4922
rect 2874 4870 2876 4922
rect 2714 4868 2738 4870
rect 2794 4868 2818 4870
rect 2874 4868 2898 4870
rect 2658 4848 2954 4868
rect 4360 4380 4656 4400
rect 4416 4378 4440 4380
rect 4496 4378 4520 4380
rect 4576 4378 4600 4380
rect 4438 4326 4440 4378
rect 4502 4326 4514 4378
rect 4576 4326 4578 4378
rect 4416 4324 4440 4326
rect 4496 4324 4520 4326
rect 4576 4324 4600 4326
rect 4360 4304 4656 4324
rect 2658 3836 2954 3856
rect 2714 3834 2738 3836
rect 2794 3834 2818 3836
rect 2874 3834 2898 3836
rect 2736 3782 2738 3834
rect 2800 3782 2812 3834
rect 2874 3782 2876 3834
rect 2714 3780 2738 3782
rect 2794 3780 2818 3782
rect 2874 3780 2898 3782
rect 2658 3760 2954 3780
rect 4360 3292 4656 3312
rect 4416 3290 4440 3292
rect 4496 3290 4520 3292
rect 4576 3290 4600 3292
rect 4438 3238 4440 3290
rect 4502 3238 4514 3290
rect 4576 3238 4578 3290
rect 4416 3236 4440 3238
rect 4496 3236 4520 3238
rect 4576 3236 4600 3238
rect 4360 3216 4656 3236
rect 2658 2748 2954 2768
rect 2714 2746 2738 2748
rect 2794 2746 2818 2748
rect 2874 2746 2898 2748
rect 2736 2694 2738 2746
rect 2800 2694 2812 2746
rect 2874 2694 2876 2746
rect 2714 2692 2738 2694
rect 2794 2692 2818 2694
rect 2874 2692 2898 2694
rect 2658 2672 2954 2692
rect 4908 2446 4936 6258
rect 6062 6012 6358 6032
rect 6118 6010 6142 6012
rect 6198 6010 6222 6012
rect 6278 6010 6302 6012
rect 6140 5958 6142 6010
rect 6204 5958 6216 6010
rect 6278 5958 6280 6010
rect 6118 5956 6142 5958
rect 6198 5956 6222 5958
rect 6278 5956 6302 5958
rect 6062 5936 6358 5956
rect 6062 4924 6358 4944
rect 6118 4922 6142 4924
rect 6198 4922 6222 4924
rect 6278 4922 6302 4924
rect 6140 4870 6142 4922
rect 6204 4870 6216 4922
rect 6278 4870 6280 4922
rect 6118 4868 6142 4870
rect 6198 4868 6222 4870
rect 6278 4868 6302 4870
rect 6062 4848 6358 4868
rect 6062 3836 6358 3856
rect 6118 3834 6142 3836
rect 6198 3834 6222 3836
rect 6278 3834 6302 3836
rect 6140 3782 6142 3834
rect 6204 3782 6216 3834
rect 6278 3782 6280 3834
rect 6118 3780 6142 3782
rect 6198 3780 6222 3782
rect 6278 3780 6302 3782
rect 6062 3760 6358 3780
rect 6062 2748 6358 2768
rect 6118 2746 6142 2748
rect 6198 2746 6222 2748
rect 6278 2746 6302 2748
rect 6140 2694 6142 2746
rect 6204 2694 6216 2746
rect 6278 2694 6280 2746
rect 6118 2692 6142 2694
rect 6198 2692 6222 2694
rect 6278 2692 6302 2694
rect 6062 2672 6358 2692
rect 7208 2446 7236 7346
rect 8956 7002 8984 7686
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9140 6798 9168 7754
rect 9466 7100 9762 7120
rect 9522 7098 9546 7100
rect 9602 7098 9626 7100
rect 9682 7098 9706 7100
rect 9544 7046 9546 7098
rect 9608 7046 9620 7098
rect 9682 7046 9684 7098
rect 9522 7044 9546 7046
rect 9602 7044 9626 7046
rect 9682 7044 9706 7046
rect 9466 7024 9762 7044
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 7764 6556 8060 6576
rect 7820 6554 7844 6556
rect 7900 6554 7924 6556
rect 7980 6554 8004 6556
rect 7842 6502 7844 6554
rect 7906 6502 7918 6554
rect 7980 6502 7982 6554
rect 7820 6500 7844 6502
rect 7900 6500 7924 6502
rect 7980 6500 8004 6502
rect 7764 6480 8060 6500
rect 9466 6012 9762 6032
rect 9522 6010 9546 6012
rect 9602 6010 9626 6012
rect 9682 6010 9706 6012
rect 9544 5958 9546 6010
rect 9608 5958 9620 6010
rect 9682 5958 9684 6010
rect 9522 5956 9546 5958
rect 9602 5956 9626 5958
rect 9682 5956 9706 5958
rect 9466 5936 9762 5956
rect 7764 5468 8060 5488
rect 7820 5466 7844 5468
rect 7900 5466 7924 5468
rect 7980 5466 8004 5468
rect 7842 5414 7844 5466
rect 7906 5414 7918 5466
rect 7980 5414 7982 5466
rect 7820 5412 7844 5414
rect 7900 5412 7924 5414
rect 7980 5412 8004 5414
rect 7764 5392 8060 5412
rect 9466 4924 9762 4944
rect 9522 4922 9546 4924
rect 9602 4922 9626 4924
rect 9682 4922 9706 4924
rect 9544 4870 9546 4922
rect 9608 4870 9620 4922
rect 9682 4870 9684 4922
rect 9522 4868 9546 4870
rect 9602 4868 9626 4870
rect 9682 4868 9706 4870
rect 9466 4848 9762 4868
rect 7764 4380 8060 4400
rect 7820 4378 7844 4380
rect 7900 4378 7924 4380
rect 7980 4378 8004 4380
rect 7842 4326 7844 4378
rect 7906 4326 7918 4378
rect 7980 4326 7982 4378
rect 7820 4324 7844 4326
rect 7900 4324 7924 4326
rect 7980 4324 8004 4326
rect 7764 4304 8060 4324
rect 9466 3836 9762 3856
rect 9522 3834 9546 3836
rect 9602 3834 9626 3836
rect 9682 3834 9706 3836
rect 9544 3782 9546 3834
rect 9608 3782 9620 3834
rect 9682 3782 9684 3834
rect 9522 3780 9546 3782
rect 9602 3780 9626 3782
rect 9682 3780 9706 3782
rect 9466 3760 9762 3780
rect 7764 3292 8060 3312
rect 7820 3290 7844 3292
rect 7900 3290 7924 3292
rect 7980 3290 8004 3292
rect 7842 3238 7844 3290
rect 7906 3238 7918 3290
rect 7980 3238 7982 3290
rect 7820 3236 7844 3238
rect 7900 3236 7924 3238
rect 7980 3236 8004 3238
rect 7764 3216 8060 3236
rect 9466 2748 9762 2768
rect 9522 2746 9546 2748
rect 9602 2746 9626 2748
rect 9682 2746 9706 2748
rect 9544 2694 9546 2746
rect 9608 2694 9620 2746
rect 9682 2694 9684 2746
rect 9522 2692 9546 2694
rect 9602 2692 9626 2694
rect 9682 2692 9706 2694
rect 9466 2672 9762 2692
rect 10336 2582 10364 7890
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 6276 2372 6328 2378
rect 6276 2314 6328 2320
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 32 800 60 2314
rect 4360 2204 4656 2224
rect 4416 2202 4440 2204
rect 4496 2202 4520 2204
rect 4576 2202 4600 2204
rect 4438 2150 4440 2202
rect 4502 2150 4514 2202
rect 4576 2150 4578 2202
rect 4416 2148 4440 2150
rect 4496 2148 4520 2150
rect 4576 2148 4600 2150
rect 4360 2128 4656 2148
rect 6288 800 6316 2314
rect 7764 2204 8060 2224
rect 7820 2202 7844 2204
rect 7900 2202 7924 2204
rect 7980 2202 8004 2204
rect 7842 2150 7844 2202
rect 7906 2150 7918 2202
rect 7980 2150 7982 2202
rect 7820 2148 7844 2150
rect 7900 2148 7924 2150
rect 7980 2148 8004 2150
rect 7764 2128 8060 2148
rect 18 0 74 800
rect 6274 0 6330 800
rect 10520 377 10548 2314
rect 10506 368 10562 377
rect 10506 303 10562 312
<< via2 >>
rect 4360 11994 4416 11996
rect 4440 11994 4496 11996
rect 4520 11994 4576 11996
rect 4600 11994 4656 11996
rect 4360 11942 4386 11994
rect 4386 11942 4416 11994
rect 4440 11942 4450 11994
rect 4450 11942 4496 11994
rect 4520 11942 4566 11994
rect 4566 11942 4576 11994
rect 4600 11942 4630 11994
rect 4630 11942 4656 11994
rect 4360 11940 4416 11942
rect 4440 11940 4496 11942
rect 4520 11940 4576 11942
rect 4600 11940 4656 11942
rect 7764 11994 7820 11996
rect 7844 11994 7900 11996
rect 7924 11994 7980 11996
rect 8004 11994 8060 11996
rect 7764 11942 7790 11994
rect 7790 11942 7820 11994
rect 7844 11942 7854 11994
rect 7854 11942 7900 11994
rect 7924 11942 7970 11994
rect 7970 11942 7980 11994
rect 8004 11942 8034 11994
rect 8034 11942 8060 11994
rect 7764 11940 7820 11942
rect 7844 11940 7900 11942
rect 7924 11940 7980 11942
rect 8004 11940 8060 11942
rect 2658 11450 2714 11452
rect 2738 11450 2794 11452
rect 2818 11450 2874 11452
rect 2898 11450 2954 11452
rect 2658 11398 2684 11450
rect 2684 11398 2714 11450
rect 2738 11398 2748 11450
rect 2748 11398 2794 11450
rect 2818 11398 2864 11450
rect 2864 11398 2874 11450
rect 2898 11398 2928 11450
rect 2928 11398 2954 11450
rect 2658 11396 2714 11398
rect 2738 11396 2794 11398
rect 2818 11396 2874 11398
rect 2898 11396 2954 11398
rect 2658 10362 2714 10364
rect 2738 10362 2794 10364
rect 2818 10362 2874 10364
rect 2898 10362 2954 10364
rect 2658 10310 2684 10362
rect 2684 10310 2714 10362
rect 2738 10310 2748 10362
rect 2748 10310 2794 10362
rect 2818 10310 2864 10362
rect 2864 10310 2874 10362
rect 2898 10310 2928 10362
rect 2928 10310 2954 10362
rect 2658 10308 2714 10310
rect 2738 10308 2794 10310
rect 2818 10308 2874 10310
rect 2898 10308 2954 10310
rect 1858 9324 1860 9344
rect 1860 9324 1912 9344
rect 1912 9324 1914 9344
rect 1858 9288 1914 9324
rect 2658 9274 2714 9276
rect 2738 9274 2794 9276
rect 2818 9274 2874 9276
rect 2898 9274 2954 9276
rect 2658 9222 2684 9274
rect 2684 9222 2714 9274
rect 2738 9222 2748 9274
rect 2748 9222 2794 9274
rect 2818 9222 2864 9274
rect 2864 9222 2874 9274
rect 2898 9222 2928 9274
rect 2928 9222 2954 9274
rect 2658 9220 2714 9222
rect 2738 9220 2794 9222
rect 2818 9220 2874 9222
rect 2898 9220 2954 9222
rect 6062 11450 6118 11452
rect 6142 11450 6198 11452
rect 6222 11450 6278 11452
rect 6302 11450 6358 11452
rect 6062 11398 6088 11450
rect 6088 11398 6118 11450
rect 6142 11398 6152 11450
rect 6152 11398 6198 11450
rect 6222 11398 6268 11450
rect 6268 11398 6278 11450
rect 6302 11398 6332 11450
rect 6332 11398 6358 11450
rect 6062 11396 6118 11398
rect 6142 11396 6198 11398
rect 6222 11396 6278 11398
rect 6302 11396 6358 11398
rect 4360 10906 4416 10908
rect 4440 10906 4496 10908
rect 4520 10906 4576 10908
rect 4600 10906 4656 10908
rect 4360 10854 4386 10906
rect 4386 10854 4416 10906
rect 4440 10854 4450 10906
rect 4450 10854 4496 10906
rect 4520 10854 4566 10906
rect 4566 10854 4576 10906
rect 4600 10854 4630 10906
rect 4630 10854 4656 10906
rect 4360 10852 4416 10854
rect 4440 10852 4496 10854
rect 4520 10852 4576 10854
rect 4600 10852 4656 10854
rect 7764 10906 7820 10908
rect 7844 10906 7900 10908
rect 7924 10906 7980 10908
rect 8004 10906 8060 10908
rect 7764 10854 7790 10906
rect 7790 10854 7820 10906
rect 7844 10854 7854 10906
rect 7854 10854 7900 10906
rect 7924 10854 7970 10906
rect 7970 10854 7980 10906
rect 8004 10854 8034 10906
rect 8034 10854 8060 10906
rect 7764 10852 7820 10854
rect 7844 10852 7900 10854
rect 7924 10852 7980 10854
rect 8004 10852 8060 10854
rect 6062 10362 6118 10364
rect 6142 10362 6198 10364
rect 6222 10362 6278 10364
rect 6302 10362 6358 10364
rect 6062 10310 6088 10362
rect 6088 10310 6118 10362
rect 6142 10310 6152 10362
rect 6152 10310 6198 10362
rect 6222 10310 6268 10362
rect 6268 10310 6278 10362
rect 6302 10310 6332 10362
rect 6332 10310 6358 10362
rect 6062 10308 6118 10310
rect 6142 10308 6198 10310
rect 6222 10308 6278 10310
rect 6302 10308 6358 10310
rect 9466 11450 9522 11452
rect 9546 11450 9602 11452
rect 9626 11450 9682 11452
rect 9706 11450 9762 11452
rect 9466 11398 9492 11450
rect 9492 11398 9522 11450
rect 9546 11398 9556 11450
rect 9556 11398 9602 11450
rect 9626 11398 9672 11450
rect 9672 11398 9682 11450
rect 9706 11398 9736 11450
rect 9736 11398 9762 11450
rect 9466 11396 9522 11398
rect 9546 11396 9602 11398
rect 9626 11396 9682 11398
rect 9706 11396 9762 11398
rect 9466 10362 9522 10364
rect 9546 10362 9602 10364
rect 9626 10362 9682 10364
rect 9706 10362 9762 10364
rect 9466 10310 9492 10362
rect 9492 10310 9522 10362
rect 9546 10310 9556 10362
rect 9556 10310 9602 10362
rect 9626 10310 9672 10362
rect 9672 10310 9682 10362
rect 9706 10310 9736 10362
rect 9736 10310 9762 10362
rect 9466 10308 9522 10310
rect 9546 10308 9602 10310
rect 9626 10308 9682 10310
rect 9706 10308 9762 10310
rect 2658 8186 2714 8188
rect 2738 8186 2794 8188
rect 2818 8186 2874 8188
rect 2898 8186 2954 8188
rect 2658 8134 2684 8186
rect 2684 8134 2714 8186
rect 2738 8134 2748 8186
rect 2748 8134 2794 8186
rect 2818 8134 2864 8186
rect 2864 8134 2874 8186
rect 2898 8134 2928 8186
rect 2928 8134 2954 8186
rect 2658 8132 2714 8134
rect 2738 8132 2794 8134
rect 2818 8132 2874 8134
rect 2898 8132 2954 8134
rect 4360 9818 4416 9820
rect 4440 9818 4496 9820
rect 4520 9818 4576 9820
rect 4600 9818 4656 9820
rect 4360 9766 4386 9818
rect 4386 9766 4416 9818
rect 4440 9766 4450 9818
rect 4450 9766 4496 9818
rect 4520 9766 4566 9818
rect 4566 9766 4576 9818
rect 4600 9766 4630 9818
rect 4630 9766 4656 9818
rect 4360 9764 4416 9766
rect 4440 9764 4496 9766
rect 4520 9764 4576 9766
rect 4600 9764 4656 9766
rect 2658 7098 2714 7100
rect 2738 7098 2794 7100
rect 2818 7098 2874 7100
rect 2898 7098 2954 7100
rect 2658 7046 2684 7098
rect 2684 7046 2714 7098
rect 2738 7046 2748 7098
rect 2748 7046 2794 7098
rect 2818 7046 2864 7098
rect 2864 7046 2874 7098
rect 2898 7046 2928 7098
rect 2928 7046 2954 7098
rect 2658 7044 2714 7046
rect 2738 7044 2794 7046
rect 2818 7044 2874 7046
rect 2898 7044 2954 7046
rect 4360 8730 4416 8732
rect 4440 8730 4496 8732
rect 4520 8730 4576 8732
rect 4600 8730 4656 8732
rect 4360 8678 4386 8730
rect 4386 8678 4416 8730
rect 4440 8678 4450 8730
rect 4450 8678 4496 8730
rect 4520 8678 4566 8730
rect 4566 8678 4576 8730
rect 4600 8678 4630 8730
rect 4630 8678 4656 8730
rect 4360 8676 4416 8678
rect 4440 8676 4496 8678
rect 4520 8676 4576 8678
rect 4600 8676 4656 8678
rect 4360 7642 4416 7644
rect 4440 7642 4496 7644
rect 4520 7642 4576 7644
rect 4600 7642 4656 7644
rect 4360 7590 4386 7642
rect 4386 7590 4416 7642
rect 4440 7590 4450 7642
rect 4450 7590 4496 7642
rect 4520 7590 4566 7642
rect 4566 7590 4576 7642
rect 4600 7590 4630 7642
rect 4630 7590 4656 7642
rect 4360 7588 4416 7590
rect 4440 7588 4496 7590
rect 4520 7588 4576 7590
rect 4600 7588 4656 7590
rect 4360 6554 4416 6556
rect 4440 6554 4496 6556
rect 4520 6554 4576 6556
rect 4600 6554 4656 6556
rect 4360 6502 4386 6554
rect 4386 6502 4416 6554
rect 4440 6502 4450 6554
rect 4450 6502 4496 6554
rect 4520 6502 4566 6554
rect 4566 6502 4576 6554
rect 4600 6502 4630 6554
rect 4630 6502 4656 6554
rect 4360 6500 4416 6502
rect 4440 6500 4496 6502
rect 4520 6500 4576 6502
rect 4600 6500 4656 6502
rect 6062 9274 6118 9276
rect 6142 9274 6198 9276
rect 6222 9274 6278 9276
rect 6302 9274 6358 9276
rect 6062 9222 6088 9274
rect 6088 9222 6118 9274
rect 6142 9222 6152 9274
rect 6152 9222 6198 9274
rect 6222 9222 6268 9274
rect 6268 9222 6278 9274
rect 6302 9222 6332 9274
rect 6332 9222 6358 9274
rect 6062 9220 6118 9222
rect 6142 9220 6198 9222
rect 6222 9220 6278 9222
rect 6302 9220 6358 9222
rect 6062 8186 6118 8188
rect 6142 8186 6198 8188
rect 6222 8186 6278 8188
rect 6302 8186 6358 8188
rect 6062 8134 6088 8186
rect 6088 8134 6118 8186
rect 6142 8134 6152 8186
rect 6152 8134 6198 8186
rect 6222 8134 6268 8186
rect 6268 8134 6278 8186
rect 6302 8134 6332 8186
rect 6332 8134 6358 8186
rect 6062 8132 6118 8134
rect 6142 8132 6198 8134
rect 6222 8132 6278 8134
rect 6302 8132 6358 8134
rect 6062 7098 6118 7100
rect 6142 7098 6198 7100
rect 6222 7098 6278 7100
rect 6302 7098 6358 7100
rect 6062 7046 6088 7098
rect 6088 7046 6118 7098
rect 6142 7046 6152 7098
rect 6152 7046 6198 7098
rect 6222 7046 6268 7098
rect 6268 7046 6278 7098
rect 6302 7046 6332 7098
rect 6332 7046 6358 7098
rect 6062 7044 6118 7046
rect 6142 7044 6198 7046
rect 6222 7044 6278 7046
rect 6302 7044 6358 7046
rect 8482 9832 8538 9888
rect 7764 9818 7820 9820
rect 7844 9818 7900 9820
rect 7924 9818 7980 9820
rect 8004 9818 8060 9820
rect 7764 9766 7790 9818
rect 7790 9766 7820 9818
rect 7844 9766 7854 9818
rect 7854 9766 7900 9818
rect 7924 9766 7970 9818
rect 7970 9766 7980 9818
rect 8004 9766 8034 9818
rect 8034 9766 8060 9818
rect 7764 9764 7820 9766
rect 7844 9764 7900 9766
rect 7924 9764 7980 9766
rect 8004 9764 8060 9766
rect 9466 9274 9522 9276
rect 9546 9274 9602 9276
rect 9626 9274 9682 9276
rect 9706 9274 9762 9276
rect 9466 9222 9492 9274
rect 9492 9222 9522 9274
rect 9546 9222 9556 9274
rect 9556 9222 9602 9274
rect 9626 9222 9672 9274
rect 9672 9222 9682 9274
rect 9706 9222 9736 9274
rect 9736 9222 9762 9274
rect 9466 9220 9522 9222
rect 9546 9220 9602 9222
rect 9626 9220 9682 9222
rect 9706 9220 9762 9222
rect 7764 8730 7820 8732
rect 7844 8730 7900 8732
rect 7924 8730 7980 8732
rect 8004 8730 8060 8732
rect 7764 8678 7790 8730
rect 7790 8678 7820 8730
rect 7844 8678 7854 8730
rect 7854 8678 7900 8730
rect 7924 8678 7970 8730
rect 7970 8678 7980 8730
rect 8004 8678 8034 8730
rect 8034 8678 8060 8730
rect 7764 8676 7820 8678
rect 7844 8676 7900 8678
rect 7924 8676 7980 8678
rect 8004 8676 8060 8678
rect 7764 7642 7820 7644
rect 7844 7642 7900 7644
rect 7924 7642 7980 7644
rect 8004 7642 8060 7644
rect 7764 7590 7790 7642
rect 7790 7590 7820 7642
rect 7844 7590 7854 7642
rect 7854 7590 7900 7642
rect 7924 7590 7970 7642
rect 7970 7590 7980 7642
rect 8004 7590 8034 7642
rect 8034 7590 8060 7642
rect 7764 7588 7820 7590
rect 7844 7588 7900 7590
rect 7924 7588 7980 7590
rect 8004 7588 8060 7590
rect 9466 8186 9522 8188
rect 9546 8186 9602 8188
rect 9626 8186 9682 8188
rect 9706 8186 9762 8188
rect 9466 8134 9492 8186
rect 9492 8134 9522 8186
rect 9546 8134 9556 8186
rect 9556 8134 9602 8186
rect 9626 8134 9672 8186
rect 9672 8134 9682 8186
rect 9706 8134 9736 8186
rect 9736 8134 9762 8186
rect 9466 8132 9522 8134
rect 9546 8132 9602 8134
rect 9626 8132 9682 8134
rect 9706 8132 9762 8134
rect 2658 6010 2714 6012
rect 2738 6010 2794 6012
rect 2818 6010 2874 6012
rect 2898 6010 2954 6012
rect 2658 5958 2684 6010
rect 2684 5958 2714 6010
rect 2738 5958 2748 6010
rect 2748 5958 2794 6010
rect 2818 5958 2864 6010
rect 2864 5958 2874 6010
rect 2898 5958 2928 6010
rect 2928 5958 2954 6010
rect 2658 5956 2714 5958
rect 2738 5956 2794 5958
rect 2818 5956 2874 5958
rect 2898 5956 2954 5958
rect 4360 5466 4416 5468
rect 4440 5466 4496 5468
rect 4520 5466 4576 5468
rect 4600 5466 4656 5468
rect 4360 5414 4386 5466
rect 4386 5414 4416 5466
rect 4440 5414 4450 5466
rect 4450 5414 4496 5466
rect 4520 5414 4566 5466
rect 4566 5414 4576 5466
rect 4600 5414 4630 5466
rect 4630 5414 4656 5466
rect 4360 5412 4416 5414
rect 4440 5412 4496 5414
rect 4520 5412 4576 5414
rect 4600 5412 4656 5414
rect 2658 4922 2714 4924
rect 2738 4922 2794 4924
rect 2818 4922 2874 4924
rect 2898 4922 2954 4924
rect 2658 4870 2684 4922
rect 2684 4870 2714 4922
rect 2738 4870 2748 4922
rect 2748 4870 2794 4922
rect 2818 4870 2864 4922
rect 2864 4870 2874 4922
rect 2898 4870 2928 4922
rect 2928 4870 2954 4922
rect 2658 4868 2714 4870
rect 2738 4868 2794 4870
rect 2818 4868 2874 4870
rect 2898 4868 2954 4870
rect 4360 4378 4416 4380
rect 4440 4378 4496 4380
rect 4520 4378 4576 4380
rect 4600 4378 4656 4380
rect 4360 4326 4386 4378
rect 4386 4326 4416 4378
rect 4440 4326 4450 4378
rect 4450 4326 4496 4378
rect 4520 4326 4566 4378
rect 4566 4326 4576 4378
rect 4600 4326 4630 4378
rect 4630 4326 4656 4378
rect 4360 4324 4416 4326
rect 4440 4324 4496 4326
rect 4520 4324 4576 4326
rect 4600 4324 4656 4326
rect 2658 3834 2714 3836
rect 2738 3834 2794 3836
rect 2818 3834 2874 3836
rect 2898 3834 2954 3836
rect 2658 3782 2684 3834
rect 2684 3782 2714 3834
rect 2738 3782 2748 3834
rect 2748 3782 2794 3834
rect 2818 3782 2864 3834
rect 2864 3782 2874 3834
rect 2898 3782 2928 3834
rect 2928 3782 2954 3834
rect 2658 3780 2714 3782
rect 2738 3780 2794 3782
rect 2818 3780 2874 3782
rect 2898 3780 2954 3782
rect 4360 3290 4416 3292
rect 4440 3290 4496 3292
rect 4520 3290 4576 3292
rect 4600 3290 4656 3292
rect 4360 3238 4386 3290
rect 4386 3238 4416 3290
rect 4440 3238 4450 3290
rect 4450 3238 4496 3290
rect 4520 3238 4566 3290
rect 4566 3238 4576 3290
rect 4600 3238 4630 3290
rect 4630 3238 4656 3290
rect 4360 3236 4416 3238
rect 4440 3236 4496 3238
rect 4520 3236 4576 3238
rect 4600 3236 4656 3238
rect 2658 2746 2714 2748
rect 2738 2746 2794 2748
rect 2818 2746 2874 2748
rect 2898 2746 2954 2748
rect 2658 2694 2684 2746
rect 2684 2694 2714 2746
rect 2738 2694 2748 2746
rect 2748 2694 2794 2746
rect 2818 2694 2864 2746
rect 2864 2694 2874 2746
rect 2898 2694 2928 2746
rect 2928 2694 2954 2746
rect 2658 2692 2714 2694
rect 2738 2692 2794 2694
rect 2818 2692 2874 2694
rect 2898 2692 2954 2694
rect 6062 6010 6118 6012
rect 6142 6010 6198 6012
rect 6222 6010 6278 6012
rect 6302 6010 6358 6012
rect 6062 5958 6088 6010
rect 6088 5958 6118 6010
rect 6142 5958 6152 6010
rect 6152 5958 6198 6010
rect 6222 5958 6268 6010
rect 6268 5958 6278 6010
rect 6302 5958 6332 6010
rect 6332 5958 6358 6010
rect 6062 5956 6118 5958
rect 6142 5956 6198 5958
rect 6222 5956 6278 5958
rect 6302 5956 6358 5958
rect 6062 4922 6118 4924
rect 6142 4922 6198 4924
rect 6222 4922 6278 4924
rect 6302 4922 6358 4924
rect 6062 4870 6088 4922
rect 6088 4870 6118 4922
rect 6142 4870 6152 4922
rect 6152 4870 6198 4922
rect 6222 4870 6268 4922
rect 6268 4870 6278 4922
rect 6302 4870 6332 4922
rect 6332 4870 6358 4922
rect 6062 4868 6118 4870
rect 6142 4868 6198 4870
rect 6222 4868 6278 4870
rect 6302 4868 6358 4870
rect 6062 3834 6118 3836
rect 6142 3834 6198 3836
rect 6222 3834 6278 3836
rect 6302 3834 6358 3836
rect 6062 3782 6088 3834
rect 6088 3782 6118 3834
rect 6142 3782 6152 3834
rect 6152 3782 6198 3834
rect 6222 3782 6268 3834
rect 6268 3782 6278 3834
rect 6302 3782 6332 3834
rect 6332 3782 6358 3834
rect 6062 3780 6118 3782
rect 6142 3780 6198 3782
rect 6222 3780 6278 3782
rect 6302 3780 6358 3782
rect 6062 2746 6118 2748
rect 6142 2746 6198 2748
rect 6222 2746 6278 2748
rect 6302 2746 6358 2748
rect 6062 2694 6088 2746
rect 6088 2694 6118 2746
rect 6142 2694 6152 2746
rect 6152 2694 6198 2746
rect 6222 2694 6268 2746
rect 6268 2694 6278 2746
rect 6302 2694 6332 2746
rect 6332 2694 6358 2746
rect 6062 2692 6118 2694
rect 6142 2692 6198 2694
rect 6222 2692 6278 2694
rect 6302 2692 6358 2694
rect 9466 7098 9522 7100
rect 9546 7098 9602 7100
rect 9626 7098 9682 7100
rect 9706 7098 9762 7100
rect 9466 7046 9492 7098
rect 9492 7046 9522 7098
rect 9546 7046 9556 7098
rect 9556 7046 9602 7098
rect 9626 7046 9672 7098
rect 9672 7046 9682 7098
rect 9706 7046 9736 7098
rect 9736 7046 9762 7098
rect 9466 7044 9522 7046
rect 9546 7044 9602 7046
rect 9626 7044 9682 7046
rect 9706 7044 9762 7046
rect 7764 6554 7820 6556
rect 7844 6554 7900 6556
rect 7924 6554 7980 6556
rect 8004 6554 8060 6556
rect 7764 6502 7790 6554
rect 7790 6502 7820 6554
rect 7844 6502 7854 6554
rect 7854 6502 7900 6554
rect 7924 6502 7970 6554
rect 7970 6502 7980 6554
rect 8004 6502 8034 6554
rect 8034 6502 8060 6554
rect 7764 6500 7820 6502
rect 7844 6500 7900 6502
rect 7924 6500 7980 6502
rect 8004 6500 8060 6502
rect 9466 6010 9522 6012
rect 9546 6010 9602 6012
rect 9626 6010 9682 6012
rect 9706 6010 9762 6012
rect 9466 5958 9492 6010
rect 9492 5958 9522 6010
rect 9546 5958 9556 6010
rect 9556 5958 9602 6010
rect 9626 5958 9672 6010
rect 9672 5958 9682 6010
rect 9706 5958 9736 6010
rect 9736 5958 9762 6010
rect 9466 5956 9522 5958
rect 9546 5956 9602 5958
rect 9626 5956 9682 5958
rect 9706 5956 9762 5958
rect 7764 5466 7820 5468
rect 7844 5466 7900 5468
rect 7924 5466 7980 5468
rect 8004 5466 8060 5468
rect 7764 5414 7790 5466
rect 7790 5414 7820 5466
rect 7844 5414 7854 5466
rect 7854 5414 7900 5466
rect 7924 5414 7970 5466
rect 7970 5414 7980 5466
rect 8004 5414 8034 5466
rect 8034 5414 8060 5466
rect 7764 5412 7820 5414
rect 7844 5412 7900 5414
rect 7924 5412 7980 5414
rect 8004 5412 8060 5414
rect 9466 4922 9522 4924
rect 9546 4922 9602 4924
rect 9626 4922 9682 4924
rect 9706 4922 9762 4924
rect 9466 4870 9492 4922
rect 9492 4870 9522 4922
rect 9546 4870 9556 4922
rect 9556 4870 9602 4922
rect 9626 4870 9672 4922
rect 9672 4870 9682 4922
rect 9706 4870 9736 4922
rect 9736 4870 9762 4922
rect 9466 4868 9522 4870
rect 9546 4868 9602 4870
rect 9626 4868 9682 4870
rect 9706 4868 9762 4870
rect 7764 4378 7820 4380
rect 7844 4378 7900 4380
rect 7924 4378 7980 4380
rect 8004 4378 8060 4380
rect 7764 4326 7790 4378
rect 7790 4326 7820 4378
rect 7844 4326 7854 4378
rect 7854 4326 7900 4378
rect 7924 4326 7970 4378
rect 7970 4326 7980 4378
rect 8004 4326 8034 4378
rect 8034 4326 8060 4378
rect 7764 4324 7820 4326
rect 7844 4324 7900 4326
rect 7924 4324 7980 4326
rect 8004 4324 8060 4326
rect 9466 3834 9522 3836
rect 9546 3834 9602 3836
rect 9626 3834 9682 3836
rect 9706 3834 9762 3836
rect 9466 3782 9492 3834
rect 9492 3782 9522 3834
rect 9546 3782 9556 3834
rect 9556 3782 9602 3834
rect 9626 3782 9672 3834
rect 9672 3782 9682 3834
rect 9706 3782 9736 3834
rect 9736 3782 9762 3834
rect 9466 3780 9522 3782
rect 9546 3780 9602 3782
rect 9626 3780 9682 3782
rect 9706 3780 9762 3782
rect 7764 3290 7820 3292
rect 7844 3290 7900 3292
rect 7924 3290 7980 3292
rect 8004 3290 8060 3292
rect 7764 3238 7790 3290
rect 7790 3238 7820 3290
rect 7844 3238 7854 3290
rect 7854 3238 7900 3290
rect 7924 3238 7970 3290
rect 7970 3238 7980 3290
rect 8004 3238 8034 3290
rect 8034 3238 8060 3290
rect 7764 3236 7820 3238
rect 7844 3236 7900 3238
rect 7924 3236 7980 3238
rect 8004 3236 8060 3238
rect 9466 2746 9522 2748
rect 9546 2746 9602 2748
rect 9626 2746 9682 2748
rect 9706 2746 9762 2748
rect 9466 2694 9492 2746
rect 9492 2694 9522 2746
rect 9546 2694 9556 2746
rect 9556 2694 9602 2746
rect 9626 2694 9672 2746
rect 9672 2694 9682 2746
rect 9706 2694 9736 2746
rect 9736 2694 9762 2746
rect 9466 2692 9522 2694
rect 9546 2692 9602 2694
rect 9626 2692 9682 2694
rect 9706 2692 9762 2694
rect 4360 2202 4416 2204
rect 4440 2202 4496 2204
rect 4520 2202 4576 2204
rect 4600 2202 4656 2204
rect 4360 2150 4386 2202
rect 4386 2150 4416 2202
rect 4440 2150 4450 2202
rect 4450 2150 4496 2202
rect 4520 2150 4566 2202
rect 4566 2150 4576 2202
rect 4600 2150 4630 2202
rect 4630 2150 4656 2202
rect 4360 2148 4416 2150
rect 4440 2148 4496 2150
rect 4520 2148 4576 2150
rect 4600 2148 4656 2150
rect 7764 2202 7820 2204
rect 7844 2202 7900 2204
rect 7924 2202 7980 2204
rect 8004 2202 8060 2204
rect 7764 2150 7790 2202
rect 7790 2150 7820 2202
rect 7844 2150 7854 2202
rect 7854 2150 7900 2202
rect 7924 2150 7970 2202
rect 7970 2150 7980 2202
rect 8004 2150 8034 2202
rect 8034 2150 8060 2202
rect 7764 2148 7820 2150
rect 7844 2148 7900 2150
rect 7924 2148 7980 2150
rect 8004 2148 8060 2150
rect 10506 312 10562 368
<< metal3 >>
rect 4348 12000 4668 12001
rect 4348 11936 4356 12000
rect 4420 11936 4436 12000
rect 4500 11936 4516 12000
rect 4580 11936 4596 12000
rect 4660 11936 4668 12000
rect 4348 11935 4668 11936
rect 7752 12000 8072 12001
rect 7752 11936 7760 12000
rect 7824 11936 7840 12000
rect 7904 11936 7920 12000
rect 7984 11936 8000 12000
rect 8064 11936 8072 12000
rect 7752 11935 8072 11936
rect 2646 11456 2966 11457
rect 2646 11392 2654 11456
rect 2718 11392 2734 11456
rect 2798 11392 2814 11456
rect 2878 11392 2894 11456
rect 2958 11392 2966 11456
rect 2646 11391 2966 11392
rect 6050 11456 6370 11457
rect 6050 11392 6058 11456
rect 6122 11392 6138 11456
rect 6202 11392 6218 11456
rect 6282 11392 6298 11456
rect 6362 11392 6370 11456
rect 6050 11391 6370 11392
rect 9454 11456 9774 11457
rect 9454 11392 9462 11456
rect 9526 11392 9542 11456
rect 9606 11392 9622 11456
rect 9686 11392 9702 11456
rect 9766 11392 9774 11456
rect 9454 11391 9774 11392
rect 4348 10912 4668 10913
rect 4348 10848 4356 10912
rect 4420 10848 4436 10912
rect 4500 10848 4516 10912
rect 4580 10848 4596 10912
rect 4660 10848 4668 10912
rect 4348 10847 4668 10848
rect 7752 10912 8072 10913
rect 7752 10848 7760 10912
rect 7824 10848 7840 10912
rect 7904 10848 7920 10912
rect 7984 10848 8000 10912
rect 8064 10848 8072 10912
rect 7752 10847 8072 10848
rect 2646 10368 2966 10369
rect 2646 10304 2654 10368
rect 2718 10304 2734 10368
rect 2798 10304 2814 10368
rect 2878 10304 2894 10368
rect 2958 10304 2966 10368
rect 2646 10303 2966 10304
rect 6050 10368 6370 10369
rect 6050 10304 6058 10368
rect 6122 10304 6138 10368
rect 6202 10304 6218 10368
rect 6282 10304 6298 10368
rect 6362 10304 6370 10368
rect 6050 10303 6370 10304
rect 9454 10368 9774 10369
rect 9454 10304 9462 10368
rect 9526 10304 9542 10368
rect 9606 10304 9622 10368
rect 9686 10304 9702 10368
rect 9766 10304 9774 10368
rect 9454 10303 9774 10304
rect 8477 9890 8543 9893
rect 11635 9890 12435 9920
rect 8477 9888 12435 9890
rect 8477 9832 8482 9888
rect 8538 9832 12435 9888
rect 8477 9830 12435 9832
rect 8477 9827 8543 9830
rect 4348 9824 4668 9825
rect 4348 9760 4356 9824
rect 4420 9760 4436 9824
rect 4500 9760 4516 9824
rect 4580 9760 4596 9824
rect 4660 9760 4668 9824
rect 4348 9759 4668 9760
rect 7752 9824 8072 9825
rect 7752 9760 7760 9824
rect 7824 9760 7840 9824
rect 7904 9760 7920 9824
rect 7984 9760 8000 9824
rect 8064 9760 8072 9824
rect 11635 9800 12435 9830
rect 7752 9759 8072 9760
rect 0 9346 800 9376
rect 1853 9346 1919 9349
rect 0 9344 1919 9346
rect 0 9288 1858 9344
rect 1914 9288 1919 9344
rect 0 9286 1919 9288
rect 0 9256 800 9286
rect 1853 9283 1919 9286
rect 2646 9280 2966 9281
rect 2646 9216 2654 9280
rect 2718 9216 2734 9280
rect 2798 9216 2814 9280
rect 2878 9216 2894 9280
rect 2958 9216 2966 9280
rect 2646 9215 2966 9216
rect 6050 9280 6370 9281
rect 6050 9216 6058 9280
rect 6122 9216 6138 9280
rect 6202 9216 6218 9280
rect 6282 9216 6298 9280
rect 6362 9216 6370 9280
rect 6050 9215 6370 9216
rect 9454 9280 9774 9281
rect 9454 9216 9462 9280
rect 9526 9216 9542 9280
rect 9606 9216 9622 9280
rect 9686 9216 9702 9280
rect 9766 9216 9774 9280
rect 9454 9215 9774 9216
rect 4348 8736 4668 8737
rect 4348 8672 4356 8736
rect 4420 8672 4436 8736
rect 4500 8672 4516 8736
rect 4580 8672 4596 8736
rect 4660 8672 4668 8736
rect 4348 8671 4668 8672
rect 7752 8736 8072 8737
rect 7752 8672 7760 8736
rect 7824 8672 7840 8736
rect 7904 8672 7920 8736
rect 7984 8672 8000 8736
rect 8064 8672 8072 8736
rect 7752 8671 8072 8672
rect 2646 8192 2966 8193
rect 2646 8128 2654 8192
rect 2718 8128 2734 8192
rect 2798 8128 2814 8192
rect 2878 8128 2894 8192
rect 2958 8128 2966 8192
rect 2646 8127 2966 8128
rect 6050 8192 6370 8193
rect 6050 8128 6058 8192
rect 6122 8128 6138 8192
rect 6202 8128 6218 8192
rect 6282 8128 6298 8192
rect 6362 8128 6370 8192
rect 6050 8127 6370 8128
rect 9454 8192 9774 8193
rect 9454 8128 9462 8192
rect 9526 8128 9542 8192
rect 9606 8128 9622 8192
rect 9686 8128 9702 8192
rect 9766 8128 9774 8192
rect 9454 8127 9774 8128
rect 4348 7648 4668 7649
rect 4348 7584 4356 7648
rect 4420 7584 4436 7648
rect 4500 7584 4516 7648
rect 4580 7584 4596 7648
rect 4660 7584 4668 7648
rect 4348 7583 4668 7584
rect 7752 7648 8072 7649
rect 7752 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8072 7648
rect 7752 7583 8072 7584
rect 2646 7104 2966 7105
rect 2646 7040 2654 7104
rect 2718 7040 2734 7104
rect 2798 7040 2814 7104
rect 2878 7040 2894 7104
rect 2958 7040 2966 7104
rect 2646 7039 2966 7040
rect 6050 7104 6370 7105
rect 6050 7040 6058 7104
rect 6122 7040 6138 7104
rect 6202 7040 6218 7104
rect 6282 7040 6298 7104
rect 6362 7040 6370 7104
rect 6050 7039 6370 7040
rect 9454 7104 9774 7105
rect 9454 7040 9462 7104
rect 9526 7040 9542 7104
rect 9606 7040 9622 7104
rect 9686 7040 9702 7104
rect 9766 7040 9774 7104
rect 9454 7039 9774 7040
rect 4348 6560 4668 6561
rect 4348 6496 4356 6560
rect 4420 6496 4436 6560
rect 4500 6496 4516 6560
rect 4580 6496 4596 6560
rect 4660 6496 4668 6560
rect 4348 6495 4668 6496
rect 7752 6560 8072 6561
rect 7752 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8072 6560
rect 7752 6495 8072 6496
rect 2646 6016 2966 6017
rect 2646 5952 2654 6016
rect 2718 5952 2734 6016
rect 2798 5952 2814 6016
rect 2878 5952 2894 6016
rect 2958 5952 2966 6016
rect 2646 5951 2966 5952
rect 6050 6016 6370 6017
rect 6050 5952 6058 6016
rect 6122 5952 6138 6016
rect 6202 5952 6218 6016
rect 6282 5952 6298 6016
rect 6362 5952 6370 6016
rect 6050 5951 6370 5952
rect 9454 6016 9774 6017
rect 9454 5952 9462 6016
rect 9526 5952 9542 6016
rect 9606 5952 9622 6016
rect 9686 5952 9702 6016
rect 9766 5952 9774 6016
rect 9454 5951 9774 5952
rect 4348 5472 4668 5473
rect 4348 5408 4356 5472
rect 4420 5408 4436 5472
rect 4500 5408 4516 5472
rect 4580 5408 4596 5472
rect 4660 5408 4668 5472
rect 4348 5407 4668 5408
rect 7752 5472 8072 5473
rect 7752 5408 7760 5472
rect 7824 5408 7840 5472
rect 7904 5408 7920 5472
rect 7984 5408 8000 5472
rect 8064 5408 8072 5472
rect 7752 5407 8072 5408
rect 2646 4928 2966 4929
rect 2646 4864 2654 4928
rect 2718 4864 2734 4928
rect 2798 4864 2814 4928
rect 2878 4864 2894 4928
rect 2958 4864 2966 4928
rect 2646 4863 2966 4864
rect 6050 4928 6370 4929
rect 6050 4864 6058 4928
rect 6122 4864 6138 4928
rect 6202 4864 6218 4928
rect 6282 4864 6298 4928
rect 6362 4864 6370 4928
rect 6050 4863 6370 4864
rect 9454 4928 9774 4929
rect 9454 4864 9462 4928
rect 9526 4864 9542 4928
rect 9606 4864 9622 4928
rect 9686 4864 9702 4928
rect 9766 4864 9774 4928
rect 9454 4863 9774 4864
rect 4348 4384 4668 4385
rect 4348 4320 4356 4384
rect 4420 4320 4436 4384
rect 4500 4320 4516 4384
rect 4580 4320 4596 4384
rect 4660 4320 4668 4384
rect 4348 4319 4668 4320
rect 7752 4384 8072 4385
rect 7752 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8072 4384
rect 7752 4319 8072 4320
rect 2646 3840 2966 3841
rect 2646 3776 2654 3840
rect 2718 3776 2734 3840
rect 2798 3776 2814 3840
rect 2878 3776 2894 3840
rect 2958 3776 2966 3840
rect 2646 3775 2966 3776
rect 6050 3840 6370 3841
rect 6050 3776 6058 3840
rect 6122 3776 6138 3840
rect 6202 3776 6218 3840
rect 6282 3776 6298 3840
rect 6362 3776 6370 3840
rect 6050 3775 6370 3776
rect 9454 3840 9774 3841
rect 9454 3776 9462 3840
rect 9526 3776 9542 3840
rect 9606 3776 9622 3840
rect 9686 3776 9702 3840
rect 9766 3776 9774 3840
rect 9454 3775 9774 3776
rect 4348 3296 4668 3297
rect 4348 3232 4356 3296
rect 4420 3232 4436 3296
rect 4500 3232 4516 3296
rect 4580 3232 4596 3296
rect 4660 3232 4668 3296
rect 4348 3231 4668 3232
rect 7752 3296 8072 3297
rect 7752 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8072 3296
rect 7752 3231 8072 3232
rect 2646 2752 2966 2753
rect 2646 2688 2654 2752
rect 2718 2688 2734 2752
rect 2798 2688 2814 2752
rect 2878 2688 2894 2752
rect 2958 2688 2966 2752
rect 2646 2687 2966 2688
rect 6050 2752 6370 2753
rect 6050 2688 6058 2752
rect 6122 2688 6138 2752
rect 6202 2688 6218 2752
rect 6282 2688 6298 2752
rect 6362 2688 6370 2752
rect 6050 2687 6370 2688
rect 9454 2752 9774 2753
rect 9454 2688 9462 2752
rect 9526 2688 9542 2752
rect 9606 2688 9622 2752
rect 9686 2688 9702 2752
rect 9766 2688 9774 2752
rect 9454 2687 9774 2688
rect 4348 2208 4668 2209
rect 4348 2144 4356 2208
rect 4420 2144 4436 2208
rect 4500 2144 4516 2208
rect 4580 2144 4596 2208
rect 4660 2144 4668 2208
rect 4348 2143 4668 2144
rect 7752 2208 8072 2209
rect 7752 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8072 2208
rect 7752 2143 8072 2144
rect 10501 370 10567 373
rect 11635 370 12435 400
rect 10501 368 12435 370
rect 10501 312 10506 368
rect 10562 312 12435 368
rect 10501 310 12435 312
rect 10501 307 10567 310
rect 11635 280 12435 310
<< via3 >>
rect 4356 11996 4420 12000
rect 4356 11940 4360 11996
rect 4360 11940 4416 11996
rect 4416 11940 4420 11996
rect 4356 11936 4420 11940
rect 4436 11996 4500 12000
rect 4436 11940 4440 11996
rect 4440 11940 4496 11996
rect 4496 11940 4500 11996
rect 4436 11936 4500 11940
rect 4516 11996 4580 12000
rect 4516 11940 4520 11996
rect 4520 11940 4576 11996
rect 4576 11940 4580 11996
rect 4516 11936 4580 11940
rect 4596 11996 4660 12000
rect 4596 11940 4600 11996
rect 4600 11940 4656 11996
rect 4656 11940 4660 11996
rect 4596 11936 4660 11940
rect 7760 11996 7824 12000
rect 7760 11940 7764 11996
rect 7764 11940 7820 11996
rect 7820 11940 7824 11996
rect 7760 11936 7824 11940
rect 7840 11996 7904 12000
rect 7840 11940 7844 11996
rect 7844 11940 7900 11996
rect 7900 11940 7904 11996
rect 7840 11936 7904 11940
rect 7920 11996 7984 12000
rect 7920 11940 7924 11996
rect 7924 11940 7980 11996
rect 7980 11940 7984 11996
rect 7920 11936 7984 11940
rect 8000 11996 8064 12000
rect 8000 11940 8004 11996
rect 8004 11940 8060 11996
rect 8060 11940 8064 11996
rect 8000 11936 8064 11940
rect 2654 11452 2718 11456
rect 2654 11396 2658 11452
rect 2658 11396 2714 11452
rect 2714 11396 2718 11452
rect 2654 11392 2718 11396
rect 2734 11452 2798 11456
rect 2734 11396 2738 11452
rect 2738 11396 2794 11452
rect 2794 11396 2798 11452
rect 2734 11392 2798 11396
rect 2814 11452 2878 11456
rect 2814 11396 2818 11452
rect 2818 11396 2874 11452
rect 2874 11396 2878 11452
rect 2814 11392 2878 11396
rect 2894 11452 2958 11456
rect 2894 11396 2898 11452
rect 2898 11396 2954 11452
rect 2954 11396 2958 11452
rect 2894 11392 2958 11396
rect 6058 11452 6122 11456
rect 6058 11396 6062 11452
rect 6062 11396 6118 11452
rect 6118 11396 6122 11452
rect 6058 11392 6122 11396
rect 6138 11452 6202 11456
rect 6138 11396 6142 11452
rect 6142 11396 6198 11452
rect 6198 11396 6202 11452
rect 6138 11392 6202 11396
rect 6218 11452 6282 11456
rect 6218 11396 6222 11452
rect 6222 11396 6278 11452
rect 6278 11396 6282 11452
rect 6218 11392 6282 11396
rect 6298 11452 6362 11456
rect 6298 11396 6302 11452
rect 6302 11396 6358 11452
rect 6358 11396 6362 11452
rect 6298 11392 6362 11396
rect 9462 11452 9526 11456
rect 9462 11396 9466 11452
rect 9466 11396 9522 11452
rect 9522 11396 9526 11452
rect 9462 11392 9526 11396
rect 9542 11452 9606 11456
rect 9542 11396 9546 11452
rect 9546 11396 9602 11452
rect 9602 11396 9606 11452
rect 9542 11392 9606 11396
rect 9622 11452 9686 11456
rect 9622 11396 9626 11452
rect 9626 11396 9682 11452
rect 9682 11396 9686 11452
rect 9622 11392 9686 11396
rect 9702 11452 9766 11456
rect 9702 11396 9706 11452
rect 9706 11396 9762 11452
rect 9762 11396 9766 11452
rect 9702 11392 9766 11396
rect 4356 10908 4420 10912
rect 4356 10852 4360 10908
rect 4360 10852 4416 10908
rect 4416 10852 4420 10908
rect 4356 10848 4420 10852
rect 4436 10908 4500 10912
rect 4436 10852 4440 10908
rect 4440 10852 4496 10908
rect 4496 10852 4500 10908
rect 4436 10848 4500 10852
rect 4516 10908 4580 10912
rect 4516 10852 4520 10908
rect 4520 10852 4576 10908
rect 4576 10852 4580 10908
rect 4516 10848 4580 10852
rect 4596 10908 4660 10912
rect 4596 10852 4600 10908
rect 4600 10852 4656 10908
rect 4656 10852 4660 10908
rect 4596 10848 4660 10852
rect 7760 10908 7824 10912
rect 7760 10852 7764 10908
rect 7764 10852 7820 10908
rect 7820 10852 7824 10908
rect 7760 10848 7824 10852
rect 7840 10908 7904 10912
rect 7840 10852 7844 10908
rect 7844 10852 7900 10908
rect 7900 10852 7904 10908
rect 7840 10848 7904 10852
rect 7920 10908 7984 10912
rect 7920 10852 7924 10908
rect 7924 10852 7980 10908
rect 7980 10852 7984 10908
rect 7920 10848 7984 10852
rect 8000 10908 8064 10912
rect 8000 10852 8004 10908
rect 8004 10852 8060 10908
rect 8060 10852 8064 10908
rect 8000 10848 8064 10852
rect 2654 10364 2718 10368
rect 2654 10308 2658 10364
rect 2658 10308 2714 10364
rect 2714 10308 2718 10364
rect 2654 10304 2718 10308
rect 2734 10364 2798 10368
rect 2734 10308 2738 10364
rect 2738 10308 2794 10364
rect 2794 10308 2798 10364
rect 2734 10304 2798 10308
rect 2814 10364 2878 10368
rect 2814 10308 2818 10364
rect 2818 10308 2874 10364
rect 2874 10308 2878 10364
rect 2814 10304 2878 10308
rect 2894 10364 2958 10368
rect 2894 10308 2898 10364
rect 2898 10308 2954 10364
rect 2954 10308 2958 10364
rect 2894 10304 2958 10308
rect 6058 10364 6122 10368
rect 6058 10308 6062 10364
rect 6062 10308 6118 10364
rect 6118 10308 6122 10364
rect 6058 10304 6122 10308
rect 6138 10364 6202 10368
rect 6138 10308 6142 10364
rect 6142 10308 6198 10364
rect 6198 10308 6202 10364
rect 6138 10304 6202 10308
rect 6218 10364 6282 10368
rect 6218 10308 6222 10364
rect 6222 10308 6278 10364
rect 6278 10308 6282 10364
rect 6218 10304 6282 10308
rect 6298 10364 6362 10368
rect 6298 10308 6302 10364
rect 6302 10308 6358 10364
rect 6358 10308 6362 10364
rect 6298 10304 6362 10308
rect 9462 10364 9526 10368
rect 9462 10308 9466 10364
rect 9466 10308 9522 10364
rect 9522 10308 9526 10364
rect 9462 10304 9526 10308
rect 9542 10364 9606 10368
rect 9542 10308 9546 10364
rect 9546 10308 9602 10364
rect 9602 10308 9606 10364
rect 9542 10304 9606 10308
rect 9622 10364 9686 10368
rect 9622 10308 9626 10364
rect 9626 10308 9682 10364
rect 9682 10308 9686 10364
rect 9622 10304 9686 10308
rect 9702 10364 9766 10368
rect 9702 10308 9706 10364
rect 9706 10308 9762 10364
rect 9762 10308 9766 10364
rect 9702 10304 9766 10308
rect 4356 9820 4420 9824
rect 4356 9764 4360 9820
rect 4360 9764 4416 9820
rect 4416 9764 4420 9820
rect 4356 9760 4420 9764
rect 4436 9820 4500 9824
rect 4436 9764 4440 9820
rect 4440 9764 4496 9820
rect 4496 9764 4500 9820
rect 4436 9760 4500 9764
rect 4516 9820 4580 9824
rect 4516 9764 4520 9820
rect 4520 9764 4576 9820
rect 4576 9764 4580 9820
rect 4516 9760 4580 9764
rect 4596 9820 4660 9824
rect 4596 9764 4600 9820
rect 4600 9764 4656 9820
rect 4656 9764 4660 9820
rect 4596 9760 4660 9764
rect 7760 9820 7824 9824
rect 7760 9764 7764 9820
rect 7764 9764 7820 9820
rect 7820 9764 7824 9820
rect 7760 9760 7824 9764
rect 7840 9820 7904 9824
rect 7840 9764 7844 9820
rect 7844 9764 7900 9820
rect 7900 9764 7904 9820
rect 7840 9760 7904 9764
rect 7920 9820 7984 9824
rect 7920 9764 7924 9820
rect 7924 9764 7980 9820
rect 7980 9764 7984 9820
rect 7920 9760 7984 9764
rect 8000 9820 8064 9824
rect 8000 9764 8004 9820
rect 8004 9764 8060 9820
rect 8060 9764 8064 9820
rect 8000 9760 8064 9764
rect 2654 9276 2718 9280
rect 2654 9220 2658 9276
rect 2658 9220 2714 9276
rect 2714 9220 2718 9276
rect 2654 9216 2718 9220
rect 2734 9276 2798 9280
rect 2734 9220 2738 9276
rect 2738 9220 2794 9276
rect 2794 9220 2798 9276
rect 2734 9216 2798 9220
rect 2814 9276 2878 9280
rect 2814 9220 2818 9276
rect 2818 9220 2874 9276
rect 2874 9220 2878 9276
rect 2814 9216 2878 9220
rect 2894 9276 2958 9280
rect 2894 9220 2898 9276
rect 2898 9220 2954 9276
rect 2954 9220 2958 9276
rect 2894 9216 2958 9220
rect 6058 9276 6122 9280
rect 6058 9220 6062 9276
rect 6062 9220 6118 9276
rect 6118 9220 6122 9276
rect 6058 9216 6122 9220
rect 6138 9276 6202 9280
rect 6138 9220 6142 9276
rect 6142 9220 6198 9276
rect 6198 9220 6202 9276
rect 6138 9216 6202 9220
rect 6218 9276 6282 9280
rect 6218 9220 6222 9276
rect 6222 9220 6278 9276
rect 6278 9220 6282 9276
rect 6218 9216 6282 9220
rect 6298 9276 6362 9280
rect 6298 9220 6302 9276
rect 6302 9220 6358 9276
rect 6358 9220 6362 9276
rect 6298 9216 6362 9220
rect 9462 9276 9526 9280
rect 9462 9220 9466 9276
rect 9466 9220 9522 9276
rect 9522 9220 9526 9276
rect 9462 9216 9526 9220
rect 9542 9276 9606 9280
rect 9542 9220 9546 9276
rect 9546 9220 9602 9276
rect 9602 9220 9606 9276
rect 9542 9216 9606 9220
rect 9622 9276 9686 9280
rect 9622 9220 9626 9276
rect 9626 9220 9682 9276
rect 9682 9220 9686 9276
rect 9622 9216 9686 9220
rect 9702 9276 9766 9280
rect 9702 9220 9706 9276
rect 9706 9220 9762 9276
rect 9762 9220 9766 9276
rect 9702 9216 9766 9220
rect 4356 8732 4420 8736
rect 4356 8676 4360 8732
rect 4360 8676 4416 8732
rect 4416 8676 4420 8732
rect 4356 8672 4420 8676
rect 4436 8732 4500 8736
rect 4436 8676 4440 8732
rect 4440 8676 4496 8732
rect 4496 8676 4500 8732
rect 4436 8672 4500 8676
rect 4516 8732 4580 8736
rect 4516 8676 4520 8732
rect 4520 8676 4576 8732
rect 4576 8676 4580 8732
rect 4516 8672 4580 8676
rect 4596 8732 4660 8736
rect 4596 8676 4600 8732
rect 4600 8676 4656 8732
rect 4656 8676 4660 8732
rect 4596 8672 4660 8676
rect 7760 8732 7824 8736
rect 7760 8676 7764 8732
rect 7764 8676 7820 8732
rect 7820 8676 7824 8732
rect 7760 8672 7824 8676
rect 7840 8732 7904 8736
rect 7840 8676 7844 8732
rect 7844 8676 7900 8732
rect 7900 8676 7904 8732
rect 7840 8672 7904 8676
rect 7920 8732 7984 8736
rect 7920 8676 7924 8732
rect 7924 8676 7980 8732
rect 7980 8676 7984 8732
rect 7920 8672 7984 8676
rect 8000 8732 8064 8736
rect 8000 8676 8004 8732
rect 8004 8676 8060 8732
rect 8060 8676 8064 8732
rect 8000 8672 8064 8676
rect 2654 8188 2718 8192
rect 2654 8132 2658 8188
rect 2658 8132 2714 8188
rect 2714 8132 2718 8188
rect 2654 8128 2718 8132
rect 2734 8188 2798 8192
rect 2734 8132 2738 8188
rect 2738 8132 2794 8188
rect 2794 8132 2798 8188
rect 2734 8128 2798 8132
rect 2814 8188 2878 8192
rect 2814 8132 2818 8188
rect 2818 8132 2874 8188
rect 2874 8132 2878 8188
rect 2814 8128 2878 8132
rect 2894 8188 2958 8192
rect 2894 8132 2898 8188
rect 2898 8132 2954 8188
rect 2954 8132 2958 8188
rect 2894 8128 2958 8132
rect 6058 8188 6122 8192
rect 6058 8132 6062 8188
rect 6062 8132 6118 8188
rect 6118 8132 6122 8188
rect 6058 8128 6122 8132
rect 6138 8188 6202 8192
rect 6138 8132 6142 8188
rect 6142 8132 6198 8188
rect 6198 8132 6202 8188
rect 6138 8128 6202 8132
rect 6218 8188 6282 8192
rect 6218 8132 6222 8188
rect 6222 8132 6278 8188
rect 6278 8132 6282 8188
rect 6218 8128 6282 8132
rect 6298 8188 6362 8192
rect 6298 8132 6302 8188
rect 6302 8132 6358 8188
rect 6358 8132 6362 8188
rect 6298 8128 6362 8132
rect 9462 8188 9526 8192
rect 9462 8132 9466 8188
rect 9466 8132 9522 8188
rect 9522 8132 9526 8188
rect 9462 8128 9526 8132
rect 9542 8188 9606 8192
rect 9542 8132 9546 8188
rect 9546 8132 9602 8188
rect 9602 8132 9606 8188
rect 9542 8128 9606 8132
rect 9622 8188 9686 8192
rect 9622 8132 9626 8188
rect 9626 8132 9682 8188
rect 9682 8132 9686 8188
rect 9622 8128 9686 8132
rect 9702 8188 9766 8192
rect 9702 8132 9706 8188
rect 9706 8132 9762 8188
rect 9762 8132 9766 8188
rect 9702 8128 9766 8132
rect 4356 7644 4420 7648
rect 4356 7588 4360 7644
rect 4360 7588 4416 7644
rect 4416 7588 4420 7644
rect 4356 7584 4420 7588
rect 4436 7644 4500 7648
rect 4436 7588 4440 7644
rect 4440 7588 4496 7644
rect 4496 7588 4500 7644
rect 4436 7584 4500 7588
rect 4516 7644 4580 7648
rect 4516 7588 4520 7644
rect 4520 7588 4576 7644
rect 4576 7588 4580 7644
rect 4516 7584 4580 7588
rect 4596 7644 4660 7648
rect 4596 7588 4600 7644
rect 4600 7588 4656 7644
rect 4656 7588 4660 7644
rect 4596 7584 4660 7588
rect 7760 7644 7824 7648
rect 7760 7588 7764 7644
rect 7764 7588 7820 7644
rect 7820 7588 7824 7644
rect 7760 7584 7824 7588
rect 7840 7644 7904 7648
rect 7840 7588 7844 7644
rect 7844 7588 7900 7644
rect 7900 7588 7904 7644
rect 7840 7584 7904 7588
rect 7920 7644 7984 7648
rect 7920 7588 7924 7644
rect 7924 7588 7980 7644
rect 7980 7588 7984 7644
rect 7920 7584 7984 7588
rect 8000 7644 8064 7648
rect 8000 7588 8004 7644
rect 8004 7588 8060 7644
rect 8060 7588 8064 7644
rect 8000 7584 8064 7588
rect 2654 7100 2718 7104
rect 2654 7044 2658 7100
rect 2658 7044 2714 7100
rect 2714 7044 2718 7100
rect 2654 7040 2718 7044
rect 2734 7100 2798 7104
rect 2734 7044 2738 7100
rect 2738 7044 2794 7100
rect 2794 7044 2798 7100
rect 2734 7040 2798 7044
rect 2814 7100 2878 7104
rect 2814 7044 2818 7100
rect 2818 7044 2874 7100
rect 2874 7044 2878 7100
rect 2814 7040 2878 7044
rect 2894 7100 2958 7104
rect 2894 7044 2898 7100
rect 2898 7044 2954 7100
rect 2954 7044 2958 7100
rect 2894 7040 2958 7044
rect 6058 7100 6122 7104
rect 6058 7044 6062 7100
rect 6062 7044 6118 7100
rect 6118 7044 6122 7100
rect 6058 7040 6122 7044
rect 6138 7100 6202 7104
rect 6138 7044 6142 7100
rect 6142 7044 6198 7100
rect 6198 7044 6202 7100
rect 6138 7040 6202 7044
rect 6218 7100 6282 7104
rect 6218 7044 6222 7100
rect 6222 7044 6278 7100
rect 6278 7044 6282 7100
rect 6218 7040 6282 7044
rect 6298 7100 6362 7104
rect 6298 7044 6302 7100
rect 6302 7044 6358 7100
rect 6358 7044 6362 7100
rect 6298 7040 6362 7044
rect 9462 7100 9526 7104
rect 9462 7044 9466 7100
rect 9466 7044 9522 7100
rect 9522 7044 9526 7100
rect 9462 7040 9526 7044
rect 9542 7100 9606 7104
rect 9542 7044 9546 7100
rect 9546 7044 9602 7100
rect 9602 7044 9606 7100
rect 9542 7040 9606 7044
rect 9622 7100 9686 7104
rect 9622 7044 9626 7100
rect 9626 7044 9682 7100
rect 9682 7044 9686 7100
rect 9622 7040 9686 7044
rect 9702 7100 9766 7104
rect 9702 7044 9706 7100
rect 9706 7044 9762 7100
rect 9762 7044 9766 7100
rect 9702 7040 9766 7044
rect 4356 6556 4420 6560
rect 4356 6500 4360 6556
rect 4360 6500 4416 6556
rect 4416 6500 4420 6556
rect 4356 6496 4420 6500
rect 4436 6556 4500 6560
rect 4436 6500 4440 6556
rect 4440 6500 4496 6556
rect 4496 6500 4500 6556
rect 4436 6496 4500 6500
rect 4516 6556 4580 6560
rect 4516 6500 4520 6556
rect 4520 6500 4576 6556
rect 4576 6500 4580 6556
rect 4516 6496 4580 6500
rect 4596 6556 4660 6560
rect 4596 6500 4600 6556
rect 4600 6500 4656 6556
rect 4656 6500 4660 6556
rect 4596 6496 4660 6500
rect 7760 6556 7824 6560
rect 7760 6500 7764 6556
rect 7764 6500 7820 6556
rect 7820 6500 7824 6556
rect 7760 6496 7824 6500
rect 7840 6556 7904 6560
rect 7840 6500 7844 6556
rect 7844 6500 7900 6556
rect 7900 6500 7904 6556
rect 7840 6496 7904 6500
rect 7920 6556 7984 6560
rect 7920 6500 7924 6556
rect 7924 6500 7980 6556
rect 7980 6500 7984 6556
rect 7920 6496 7984 6500
rect 8000 6556 8064 6560
rect 8000 6500 8004 6556
rect 8004 6500 8060 6556
rect 8060 6500 8064 6556
rect 8000 6496 8064 6500
rect 2654 6012 2718 6016
rect 2654 5956 2658 6012
rect 2658 5956 2714 6012
rect 2714 5956 2718 6012
rect 2654 5952 2718 5956
rect 2734 6012 2798 6016
rect 2734 5956 2738 6012
rect 2738 5956 2794 6012
rect 2794 5956 2798 6012
rect 2734 5952 2798 5956
rect 2814 6012 2878 6016
rect 2814 5956 2818 6012
rect 2818 5956 2874 6012
rect 2874 5956 2878 6012
rect 2814 5952 2878 5956
rect 2894 6012 2958 6016
rect 2894 5956 2898 6012
rect 2898 5956 2954 6012
rect 2954 5956 2958 6012
rect 2894 5952 2958 5956
rect 6058 6012 6122 6016
rect 6058 5956 6062 6012
rect 6062 5956 6118 6012
rect 6118 5956 6122 6012
rect 6058 5952 6122 5956
rect 6138 6012 6202 6016
rect 6138 5956 6142 6012
rect 6142 5956 6198 6012
rect 6198 5956 6202 6012
rect 6138 5952 6202 5956
rect 6218 6012 6282 6016
rect 6218 5956 6222 6012
rect 6222 5956 6278 6012
rect 6278 5956 6282 6012
rect 6218 5952 6282 5956
rect 6298 6012 6362 6016
rect 6298 5956 6302 6012
rect 6302 5956 6358 6012
rect 6358 5956 6362 6012
rect 6298 5952 6362 5956
rect 9462 6012 9526 6016
rect 9462 5956 9466 6012
rect 9466 5956 9522 6012
rect 9522 5956 9526 6012
rect 9462 5952 9526 5956
rect 9542 6012 9606 6016
rect 9542 5956 9546 6012
rect 9546 5956 9602 6012
rect 9602 5956 9606 6012
rect 9542 5952 9606 5956
rect 9622 6012 9686 6016
rect 9622 5956 9626 6012
rect 9626 5956 9682 6012
rect 9682 5956 9686 6012
rect 9622 5952 9686 5956
rect 9702 6012 9766 6016
rect 9702 5956 9706 6012
rect 9706 5956 9762 6012
rect 9762 5956 9766 6012
rect 9702 5952 9766 5956
rect 4356 5468 4420 5472
rect 4356 5412 4360 5468
rect 4360 5412 4416 5468
rect 4416 5412 4420 5468
rect 4356 5408 4420 5412
rect 4436 5468 4500 5472
rect 4436 5412 4440 5468
rect 4440 5412 4496 5468
rect 4496 5412 4500 5468
rect 4436 5408 4500 5412
rect 4516 5468 4580 5472
rect 4516 5412 4520 5468
rect 4520 5412 4576 5468
rect 4576 5412 4580 5468
rect 4516 5408 4580 5412
rect 4596 5468 4660 5472
rect 4596 5412 4600 5468
rect 4600 5412 4656 5468
rect 4656 5412 4660 5468
rect 4596 5408 4660 5412
rect 7760 5468 7824 5472
rect 7760 5412 7764 5468
rect 7764 5412 7820 5468
rect 7820 5412 7824 5468
rect 7760 5408 7824 5412
rect 7840 5468 7904 5472
rect 7840 5412 7844 5468
rect 7844 5412 7900 5468
rect 7900 5412 7904 5468
rect 7840 5408 7904 5412
rect 7920 5468 7984 5472
rect 7920 5412 7924 5468
rect 7924 5412 7980 5468
rect 7980 5412 7984 5468
rect 7920 5408 7984 5412
rect 8000 5468 8064 5472
rect 8000 5412 8004 5468
rect 8004 5412 8060 5468
rect 8060 5412 8064 5468
rect 8000 5408 8064 5412
rect 2654 4924 2718 4928
rect 2654 4868 2658 4924
rect 2658 4868 2714 4924
rect 2714 4868 2718 4924
rect 2654 4864 2718 4868
rect 2734 4924 2798 4928
rect 2734 4868 2738 4924
rect 2738 4868 2794 4924
rect 2794 4868 2798 4924
rect 2734 4864 2798 4868
rect 2814 4924 2878 4928
rect 2814 4868 2818 4924
rect 2818 4868 2874 4924
rect 2874 4868 2878 4924
rect 2814 4864 2878 4868
rect 2894 4924 2958 4928
rect 2894 4868 2898 4924
rect 2898 4868 2954 4924
rect 2954 4868 2958 4924
rect 2894 4864 2958 4868
rect 6058 4924 6122 4928
rect 6058 4868 6062 4924
rect 6062 4868 6118 4924
rect 6118 4868 6122 4924
rect 6058 4864 6122 4868
rect 6138 4924 6202 4928
rect 6138 4868 6142 4924
rect 6142 4868 6198 4924
rect 6198 4868 6202 4924
rect 6138 4864 6202 4868
rect 6218 4924 6282 4928
rect 6218 4868 6222 4924
rect 6222 4868 6278 4924
rect 6278 4868 6282 4924
rect 6218 4864 6282 4868
rect 6298 4924 6362 4928
rect 6298 4868 6302 4924
rect 6302 4868 6358 4924
rect 6358 4868 6362 4924
rect 6298 4864 6362 4868
rect 9462 4924 9526 4928
rect 9462 4868 9466 4924
rect 9466 4868 9522 4924
rect 9522 4868 9526 4924
rect 9462 4864 9526 4868
rect 9542 4924 9606 4928
rect 9542 4868 9546 4924
rect 9546 4868 9602 4924
rect 9602 4868 9606 4924
rect 9542 4864 9606 4868
rect 9622 4924 9686 4928
rect 9622 4868 9626 4924
rect 9626 4868 9682 4924
rect 9682 4868 9686 4924
rect 9622 4864 9686 4868
rect 9702 4924 9766 4928
rect 9702 4868 9706 4924
rect 9706 4868 9762 4924
rect 9762 4868 9766 4924
rect 9702 4864 9766 4868
rect 4356 4380 4420 4384
rect 4356 4324 4360 4380
rect 4360 4324 4416 4380
rect 4416 4324 4420 4380
rect 4356 4320 4420 4324
rect 4436 4380 4500 4384
rect 4436 4324 4440 4380
rect 4440 4324 4496 4380
rect 4496 4324 4500 4380
rect 4436 4320 4500 4324
rect 4516 4380 4580 4384
rect 4516 4324 4520 4380
rect 4520 4324 4576 4380
rect 4576 4324 4580 4380
rect 4516 4320 4580 4324
rect 4596 4380 4660 4384
rect 4596 4324 4600 4380
rect 4600 4324 4656 4380
rect 4656 4324 4660 4380
rect 4596 4320 4660 4324
rect 7760 4380 7824 4384
rect 7760 4324 7764 4380
rect 7764 4324 7820 4380
rect 7820 4324 7824 4380
rect 7760 4320 7824 4324
rect 7840 4380 7904 4384
rect 7840 4324 7844 4380
rect 7844 4324 7900 4380
rect 7900 4324 7904 4380
rect 7840 4320 7904 4324
rect 7920 4380 7984 4384
rect 7920 4324 7924 4380
rect 7924 4324 7980 4380
rect 7980 4324 7984 4380
rect 7920 4320 7984 4324
rect 8000 4380 8064 4384
rect 8000 4324 8004 4380
rect 8004 4324 8060 4380
rect 8060 4324 8064 4380
rect 8000 4320 8064 4324
rect 2654 3836 2718 3840
rect 2654 3780 2658 3836
rect 2658 3780 2714 3836
rect 2714 3780 2718 3836
rect 2654 3776 2718 3780
rect 2734 3836 2798 3840
rect 2734 3780 2738 3836
rect 2738 3780 2794 3836
rect 2794 3780 2798 3836
rect 2734 3776 2798 3780
rect 2814 3836 2878 3840
rect 2814 3780 2818 3836
rect 2818 3780 2874 3836
rect 2874 3780 2878 3836
rect 2814 3776 2878 3780
rect 2894 3836 2958 3840
rect 2894 3780 2898 3836
rect 2898 3780 2954 3836
rect 2954 3780 2958 3836
rect 2894 3776 2958 3780
rect 6058 3836 6122 3840
rect 6058 3780 6062 3836
rect 6062 3780 6118 3836
rect 6118 3780 6122 3836
rect 6058 3776 6122 3780
rect 6138 3836 6202 3840
rect 6138 3780 6142 3836
rect 6142 3780 6198 3836
rect 6198 3780 6202 3836
rect 6138 3776 6202 3780
rect 6218 3836 6282 3840
rect 6218 3780 6222 3836
rect 6222 3780 6278 3836
rect 6278 3780 6282 3836
rect 6218 3776 6282 3780
rect 6298 3836 6362 3840
rect 6298 3780 6302 3836
rect 6302 3780 6358 3836
rect 6358 3780 6362 3836
rect 6298 3776 6362 3780
rect 9462 3836 9526 3840
rect 9462 3780 9466 3836
rect 9466 3780 9522 3836
rect 9522 3780 9526 3836
rect 9462 3776 9526 3780
rect 9542 3836 9606 3840
rect 9542 3780 9546 3836
rect 9546 3780 9602 3836
rect 9602 3780 9606 3836
rect 9542 3776 9606 3780
rect 9622 3836 9686 3840
rect 9622 3780 9626 3836
rect 9626 3780 9682 3836
rect 9682 3780 9686 3836
rect 9622 3776 9686 3780
rect 9702 3836 9766 3840
rect 9702 3780 9706 3836
rect 9706 3780 9762 3836
rect 9762 3780 9766 3836
rect 9702 3776 9766 3780
rect 4356 3292 4420 3296
rect 4356 3236 4360 3292
rect 4360 3236 4416 3292
rect 4416 3236 4420 3292
rect 4356 3232 4420 3236
rect 4436 3292 4500 3296
rect 4436 3236 4440 3292
rect 4440 3236 4496 3292
rect 4496 3236 4500 3292
rect 4436 3232 4500 3236
rect 4516 3292 4580 3296
rect 4516 3236 4520 3292
rect 4520 3236 4576 3292
rect 4576 3236 4580 3292
rect 4516 3232 4580 3236
rect 4596 3292 4660 3296
rect 4596 3236 4600 3292
rect 4600 3236 4656 3292
rect 4656 3236 4660 3292
rect 4596 3232 4660 3236
rect 7760 3292 7824 3296
rect 7760 3236 7764 3292
rect 7764 3236 7820 3292
rect 7820 3236 7824 3292
rect 7760 3232 7824 3236
rect 7840 3292 7904 3296
rect 7840 3236 7844 3292
rect 7844 3236 7900 3292
rect 7900 3236 7904 3292
rect 7840 3232 7904 3236
rect 7920 3292 7984 3296
rect 7920 3236 7924 3292
rect 7924 3236 7980 3292
rect 7980 3236 7984 3292
rect 7920 3232 7984 3236
rect 8000 3292 8064 3296
rect 8000 3236 8004 3292
rect 8004 3236 8060 3292
rect 8060 3236 8064 3292
rect 8000 3232 8064 3236
rect 2654 2748 2718 2752
rect 2654 2692 2658 2748
rect 2658 2692 2714 2748
rect 2714 2692 2718 2748
rect 2654 2688 2718 2692
rect 2734 2748 2798 2752
rect 2734 2692 2738 2748
rect 2738 2692 2794 2748
rect 2794 2692 2798 2748
rect 2734 2688 2798 2692
rect 2814 2748 2878 2752
rect 2814 2692 2818 2748
rect 2818 2692 2874 2748
rect 2874 2692 2878 2748
rect 2814 2688 2878 2692
rect 2894 2748 2958 2752
rect 2894 2692 2898 2748
rect 2898 2692 2954 2748
rect 2954 2692 2958 2748
rect 2894 2688 2958 2692
rect 6058 2748 6122 2752
rect 6058 2692 6062 2748
rect 6062 2692 6118 2748
rect 6118 2692 6122 2748
rect 6058 2688 6122 2692
rect 6138 2748 6202 2752
rect 6138 2692 6142 2748
rect 6142 2692 6198 2748
rect 6198 2692 6202 2748
rect 6138 2688 6202 2692
rect 6218 2748 6282 2752
rect 6218 2692 6222 2748
rect 6222 2692 6278 2748
rect 6278 2692 6282 2748
rect 6218 2688 6282 2692
rect 6298 2748 6362 2752
rect 6298 2692 6302 2748
rect 6302 2692 6358 2748
rect 6358 2692 6362 2748
rect 6298 2688 6362 2692
rect 9462 2748 9526 2752
rect 9462 2692 9466 2748
rect 9466 2692 9522 2748
rect 9522 2692 9526 2748
rect 9462 2688 9526 2692
rect 9542 2748 9606 2752
rect 9542 2692 9546 2748
rect 9546 2692 9602 2748
rect 9602 2692 9606 2748
rect 9542 2688 9606 2692
rect 9622 2748 9686 2752
rect 9622 2692 9626 2748
rect 9626 2692 9682 2748
rect 9682 2692 9686 2748
rect 9622 2688 9686 2692
rect 9702 2748 9766 2752
rect 9702 2692 9706 2748
rect 9706 2692 9762 2748
rect 9762 2692 9766 2748
rect 9702 2688 9766 2692
rect 4356 2204 4420 2208
rect 4356 2148 4360 2204
rect 4360 2148 4416 2204
rect 4416 2148 4420 2204
rect 4356 2144 4420 2148
rect 4436 2204 4500 2208
rect 4436 2148 4440 2204
rect 4440 2148 4496 2204
rect 4496 2148 4500 2204
rect 4436 2144 4500 2148
rect 4516 2204 4580 2208
rect 4516 2148 4520 2204
rect 4520 2148 4576 2204
rect 4576 2148 4580 2204
rect 4516 2144 4580 2148
rect 4596 2204 4660 2208
rect 4596 2148 4600 2204
rect 4600 2148 4656 2204
rect 4656 2148 4660 2204
rect 4596 2144 4660 2148
rect 7760 2204 7824 2208
rect 7760 2148 7764 2204
rect 7764 2148 7820 2204
rect 7820 2148 7824 2204
rect 7760 2144 7824 2148
rect 7840 2204 7904 2208
rect 7840 2148 7844 2204
rect 7844 2148 7900 2204
rect 7900 2148 7904 2204
rect 7840 2144 7904 2148
rect 7920 2204 7984 2208
rect 7920 2148 7924 2204
rect 7924 2148 7980 2204
rect 7980 2148 7984 2204
rect 7920 2144 7984 2148
rect 8000 2204 8064 2208
rect 8000 2148 8004 2204
rect 8004 2148 8060 2204
rect 8060 2148 8064 2204
rect 8000 2144 8064 2148
<< metal4 >>
rect 2646 11456 2966 12016
rect 2646 11392 2654 11456
rect 2718 11392 2734 11456
rect 2798 11392 2814 11456
rect 2878 11392 2894 11456
rect 2958 11392 2966 11456
rect 2646 10406 2966 11392
rect 2646 10368 2688 10406
rect 2924 10368 2966 10406
rect 2646 10304 2654 10368
rect 2958 10304 2966 10368
rect 2646 10170 2688 10304
rect 2924 10170 2966 10304
rect 2646 9280 2966 10170
rect 2646 9216 2654 9280
rect 2718 9216 2734 9280
rect 2798 9216 2814 9280
rect 2878 9216 2894 9280
rect 2958 9216 2966 9280
rect 2646 8192 2966 9216
rect 2646 8128 2654 8192
rect 2718 8128 2734 8192
rect 2798 8128 2814 8192
rect 2878 8128 2894 8192
rect 2958 8128 2966 8192
rect 2646 7142 2966 8128
rect 2646 7104 2688 7142
rect 2924 7104 2966 7142
rect 2646 7040 2654 7104
rect 2958 7040 2966 7104
rect 2646 6906 2688 7040
rect 2924 6906 2966 7040
rect 2646 6016 2966 6906
rect 2646 5952 2654 6016
rect 2718 5952 2734 6016
rect 2798 5952 2814 6016
rect 2878 5952 2894 6016
rect 2958 5952 2966 6016
rect 2646 4928 2966 5952
rect 2646 4864 2654 4928
rect 2718 4864 2734 4928
rect 2798 4864 2814 4928
rect 2878 4864 2894 4928
rect 2958 4864 2966 4928
rect 2646 3878 2966 4864
rect 2646 3840 2688 3878
rect 2924 3840 2966 3878
rect 2646 3776 2654 3840
rect 2958 3776 2966 3840
rect 2646 3642 2688 3776
rect 2924 3642 2966 3776
rect 2646 2752 2966 3642
rect 2646 2688 2654 2752
rect 2718 2688 2734 2752
rect 2798 2688 2814 2752
rect 2878 2688 2894 2752
rect 2958 2688 2966 2752
rect 2646 2128 2966 2688
rect 4348 12000 4668 12016
rect 4348 11936 4356 12000
rect 4420 11936 4436 12000
rect 4500 11936 4516 12000
rect 4580 11936 4596 12000
rect 4660 11936 4668 12000
rect 4348 10912 4668 11936
rect 4348 10848 4356 10912
rect 4420 10848 4436 10912
rect 4500 10848 4516 10912
rect 4580 10848 4596 10912
rect 4660 10848 4668 10912
rect 4348 9824 4668 10848
rect 4348 9760 4356 9824
rect 4420 9760 4436 9824
rect 4500 9760 4516 9824
rect 4580 9760 4596 9824
rect 4660 9760 4668 9824
rect 4348 8774 4668 9760
rect 4348 8736 4390 8774
rect 4626 8736 4668 8774
rect 4348 8672 4356 8736
rect 4660 8672 4668 8736
rect 4348 8538 4390 8672
rect 4626 8538 4668 8672
rect 4348 7648 4668 8538
rect 4348 7584 4356 7648
rect 4420 7584 4436 7648
rect 4500 7584 4516 7648
rect 4580 7584 4596 7648
rect 4660 7584 4668 7648
rect 4348 6560 4668 7584
rect 4348 6496 4356 6560
rect 4420 6496 4436 6560
rect 4500 6496 4516 6560
rect 4580 6496 4596 6560
rect 4660 6496 4668 6560
rect 4348 5510 4668 6496
rect 4348 5472 4390 5510
rect 4626 5472 4668 5510
rect 4348 5408 4356 5472
rect 4660 5408 4668 5472
rect 4348 5274 4390 5408
rect 4626 5274 4668 5408
rect 4348 4384 4668 5274
rect 4348 4320 4356 4384
rect 4420 4320 4436 4384
rect 4500 4320 4516 4384
rect 4580 4320 4596 4384
rect 4660 4320 4668 4384
rect 4348 3296 4668 4320
rect 4348 3232 4356 3296
rect 4420 3232 4436 3296
rect 4500 3232 4516 3296
rect 4580 3232 4596 3296
rect 4660 3232 4668 3296
rect 4348 2208 4668 3232
rect 4348 2144 4356 2208
rect 4420 2144 4436 2208
rect 4500 2144 4516 2208
rect 4580 2144 4596 2208
rect 4660 2144 4668 2208
rect 4348 2128 4668 2144
rect 6050 11456 6370 12016
rect 6050 11392 6058 11456
rect 6122 11392 6138 11456
rect 6202 11392 6218 11456
rect 6282 11392 6298 11456
rect 6362 11392 6370 11456
rect 6050 10406 6370 11392
rect 6050 10368 6092 10406
rect 6328 10368 6370 10406
rect 6050 10304 6058 10368
rect 6362 10304 6370 10368
rect 6050 10170 6092 10304
rect 6328 10170 6370 10304
rect 6050 9280 6370 10170
rect 6050 9216 6058 9280
rect 6122 9216 6138 9280
rect 6202 9216 6218 9280
rect 6282 9216 6298 9280
rect 6362 9216 6370 9280
rect 6050 8192 6370 9216
rect 6050 8128 6058 8192
rect 6122 8128 6138 8192
rect 6202 8128 6218 8192
rect 6282 8128 6298 8192
rect 6362 8128 6370 8192
rect 6050 7142 6370 8128
rect 6050 7104 6092 7142
rect 6328 7104 6370 7142
rect 6050 7040 6058 7104
rect 6362 7040 6370 7104
rect 6050 6906 6092 7040
rect 6328 6906 6370 7040
rect 6050 6016 6370 6906
rect 6050 5952 6058 6016
rect 6122 5952 6138 6016
rect 6202 5952 6218 6016
rect 6282 5952 6298 6016
rect 6362 5952 6370 6016
rect 6050 4928 6370 5952
rect 6050 4864 6058 4928
rect 6122 4864 6138 4928
rect 6202 4864 6218 4928
rect 6282 4864 6298 4928
rect 6362 4864 6370 4928
rect 6050 3878 6370 4864
rect 6050 3840 6092 3878
rect 6328 3840 6370 3878
rect 6050 3776 6058 3840
rect 6362 3776 6370 3840
rect 6050 3642 6092 3776
rect 6328 3642 6370 3776
rect 6050 2752 6370 3642
rect 6050 2688 6058 2752
rect 6122 2688 6138 2752
rect 6202 2688 6218 2752
rect 6282 2688 6298 2752
rect 6362 2688 6370 2752
rect 6050 2128 6370 2688
rect 7752 12000 8072 12016
rect 7752 11936 7760 12000
rect 7824 11936 7840 12000
rect 7904 11936 7920 12000
rect 7984 11936 8000 12000
rect 8064 11936 8072 12000
rect 7752 10912 8072 11936
rect 7752 10848 7760 10912
rect 7824 10848 7840 10912
rect 7904 10848 7920 10912
rect 7984 10848 8000 10912
rect 8064 10848 8072 10912
rect 7752 9824 8072 10848
rect 7752 9760 7760 9824
rect 7824 9760 7840 9824
rect 7904 9760 7920 9824
rect 7984 9760 8000 9824
rect 8064 9760 8072 9824
rect 7752 8774 8072 9760
rect 7752 8736 7794 8774
rect 8030 8736 8072 8774
rect 7752 8672 7760 8736
rect 8064 8672 8072 8736
rect 7752 8538 7794 8672
rect 8030 8538 8072 8672
rect 7752 7648 8072 8538
rect 7752 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8072 7648
rect 7752 6560 8072 7584
rect 7752 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8072 6560
rect 7752 5510 8072 6496
rect 7752 5472 7794 5510
rect 8030 5472 8072 5510
rect 7752 5408 7760 5472
rect 8064 5408 8072 5472
rect 7752 5274 7794 5408
rect 8030 5274 8072 5408
rect 7752 4384 8072 5274
rect 7752 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8072 4384
rect 7752 3296 8072 4320
rect 7752 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8072 3296
rect 7752 2208 8072 3232
rect 7752 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8072 2208
rect 7752 2128 8072 2144
rect 9454 11456 9774 12016
rect 9454 11392 9462 11456
rect 9526 11392 9542 11456
rect 9606 11392 9622 11456
rect 9686 11392 9702 11456
rect 9766 11392 9774 11456
rect 9454 10406 9774 11392
rect 9454 10368 9496 10406
rect 9732 10368 9774 10406
rect 9454 10304 9462 10368
rect 9766 10304 9774 10368
rect 9454 10170 9496 10304
rect 9732 10170 9774 10304
rect 9454 9280 9774 10170
rect 9454 9216 9462 9280
rect 9526 9216 9542 9280
rect 9606 9216 9622 9280
rect 9686 9216 9702 9280
rect 9766 9216 9774 9280
rect 9454 8192 9774 9216
rect 9454 8128 9462 8192
rect 9526 8128 9542 8192
rect 9606 8128 9622 8192
rect 9686 8128 9702 8192
rect 9766 8128 9774 8192
rect 9454 7142 9774 8128
rect 9454 7104 9496 7142
rect 9732 7104 9774 7142
rect 9454 7040 9462 7104
rect 9766 7040 9774 7104
rect 9454 6906 9496 7040
rect 9732 6906 9774 7040
rect 9454 6016 9774 6906
rect 9454 5952 9462 6016
rect 9526 5952 9542 6016
rect 9606 5952 9622 6016
rect 9686 5952 9702 6016
rect 9766 5952 9774 6016
rect 9454 4928 9774 5952
rect 9454 4864 9462 4928
rect 9526 4864 9542 4928
rect 9606 4864 9622 4928
rect 9686 4864 9702 4928
rect 9766 4864 9774 4928
rect 9454 3878 9774 4864
rect 9454 3840 9496 3878
rect 9732 3840 9774 3878
rect 9454 3776 9462 3840
rect 9766 3776 9774 3840
rect 9454 3642 9496 3776
rect 9732 3642 9774 3776
rect 9454 2752 9774 3642
rect 9454 2688 9462 2752
rect 9526 2688 9542 2752
rect 9606 2688 9622 2752
rect 9686 2688 9702 2752
rect 9766 2688 9774 2752
rect 9454 2128 9774 2688
<< via4 >>
rect 2688 10368 2924 10406
rect 2688 10304 2718 10368
rect 2718 10304 2734 10368
rect 2734 10304 2798 10368
rect 2798 10304 2814 10368
rect 2814 10304 2878 10368
rect 2878 10304 2894 10368
rect 2894 10304 2924 10368
rect 2688 10170 2924 10304
rect 2688 7104 2924 7142
rect 2688 7040 2718 7104
rect 2718 7040 2734 7104
rect 2734 7040 2798 7104
rect 2798 7040 2814 7104
rect 2814 7040 2878 7104
rect 2878 7040 2894 7104
rect 2894 7040 2924 7104
rect 2688 6906 2924 7040
rect 2688 3840 2924 3878
rect 2688 3776 2718 3840
rect 2718 3776 2734 3840
rect 2734 3776 2798 3840
rect 2798 3776 2814 3840
rect 2814 3776 2878 3840
rect 2878 3776 2894 3840
rect 2894 3776 2924 3840
rect 2688 3642 2924 3776
rect 4390 8736 4626 8774
rect 4390 8672 4420 8736
rect 4420 8672 4436 8736
rect 4436 8672 4500 8736
rect 4500 8672 4516 8736
rect 4516 8672 4580 8736
rect 4580 8672 4596 8736
rect 4596 8672 4626 8736
rect 4390 8538 4626 8672
rect 4390 5472 4626 5510
rect 4390 5408 4420 5472
rect 4420 5408 4436 5472
rect 4436 5408 4500 5472
rect 4500 5408 4516 5472
rect 4516 5408 4580 5472
rect 4580 5408 4596 5472
rect 4596 5408 4626 5472
rect 4390 5274 4626 5408
rect 6092 10368 6328 10406
rect 6092 10304 6122 10368
rect 6122 10304 6138 10368
rect 6138 10304 6202 10368
rect 6202 10304 6218 10368
rect 6218 10304 6282 10368
rect 6282 10304 6298 10368
rect 6298 10304 6328 10368
rect 6092 10170 6328 10304
rect 6092 7104 6328 7142
rect 6092 7040 6122 7104
rect 6122 7040 6138 7104
rect 6138 7040 6202 7104
rect 6202 7040 6218 7104
rect 6218 7040 6282 7104
rect 6282 7040 6298 7104
rect 6298 7040 6328 7104
rect 6092 6906 6328 7040
rect 6092 3840 6328 3878
rect 6092 3776 6122 3840
rect 6122 3776 6138 3840
rect 6138 3776 6202 3840
rect 6202 3776 6218 3840
rect 6218 3776 6282 3840
rect 6282 3776 6298 3840
rect 6298 3776 6328 3840
rect 6092 3642 6328 3776
rect 7794 8736 8030 8774
rect 7794 8672 7824 8736
rect 7824 8672 7840 8736
rect 7840 8672 7904 8736
rect 7904 8672 7920 8736
rect 7920 8672 7984 8736
rect 7984 8672 8000 8736
rect 8000 8672 8030 8736
rect 7794 8538 8030 8672
rect 7794 5472 8030 5510
rect 7794 5408 7824 5472
rect 7824 5408 7840 5472
rect 7840 5408 7904 5472
rect 7904 5408 7920 5472
rect 7920 5408 7984 5472
rect 7984 5408 8000 5472
rect 8000 5408 8030 5472
rect 7794 5274 8030 5408
rect 9496 10368 9732 10406
rect 9496 10304 9526 10368
rect 9526 10304 9542 10368
rect 9542 10304 9606 10368
rect 9606 10304 9622 10368
rect 9622 10304 9686 10368
rect 9686 10304 9702 10368
rect 9702 10304 9732 10368
rect 9496 10170 9732 10304
rect 9496 7104 9732 7142
rect 9496 7040 9526 7104
rect 9526 7040 9542 7104
rect 9542 7040 9606 7104
rect 9606 7040 9622 7104
rect 9622 7040 9686 7104
rect 9686 7040 9702 7104
rect 9702 7040 9732 7104
rect 9496 6906 9732 7040
rect 9496 3840 9732 3878
rect 9496 3776 9526 3840
rect 9526 3776 9542 3840
rect 9542 3776 9606 3840
rect 9606 3776 9622 3840
rect 9622 3776 9686 3840
rect 9686 3776 9702 3840
rect 9702 3776 9732 3840
rect 9496 3642 9732 3776
<< metal5 >>
rect 1104 10406 11316 10448
rect 1104 10170 2688 10406
rect 2924 10170 6092 10406
rect 6328 10170 9496 10406
rect 9732 10170 11316 10406
rect 1104 10128 11316 10170
rect 1104 8774 11316 8816
rect 1104 8538 4390 8774
rect 4626 8538 7794 8774
rect 8030 8538 11316 8774
rect 1104 8496 11316 8538
rect 1104 7142 11316 7184
rect 1104 6906 2688 7142
rect 2924 6906 6092 7142
rect 6328 6906 9496 7142
rect 9732 6906 11316 7142
rect 1104 6864 11316 6906
rect 1104 5510 11316 5552
rect 1104 5274 4390 5510
rect 4626 5274 7794 5510
rect 8030 5274 11316 5510
rect 1104 5232 11316 5274
rect 1104 3878 11316 3920
rect 1104 3642 2688 3878
rect 2924 3642 6092 3878
rect 6328 3642 9496 3878
rect 9732 3642 11316 3878
rect 1104 3600 11316 3642
use sky130_fd_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1629394407
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1629394407
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1629394407
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1629394407
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1629394407
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1629394407
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1629394407
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1629394407
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1629394407
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1629394407
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1629394407
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1629394407
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1629394407
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1629394407
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1629394407
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1629394407
transform -1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_65
timestamp 1629394407
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1629394407
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1629394407
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1629394407
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1629394407
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1629394407
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 1629394407
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1629394407
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1629394407
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1629394407
transform -1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp 1629394407
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1629394407
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1629394407
transform -1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1629394407
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1629394407
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1629394407
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1629394407
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1629394407
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1629394407
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1629394407
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1629394407
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1629394407
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1629394407
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1629394407
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1629394407
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1629394407
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_105
timestamp 1629394407
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1629394407
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1629394407
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1629394407
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1629394407
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1629394407
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1629394407
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1629394407
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1629394407
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1629394407
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1629394407
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1629394407
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1629394407
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1629394407
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp 1629394407
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1629394407
transform -1 0 11316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1629394407
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1629394407
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1629394407
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1629394407
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1629394407
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1629394407
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1629394407
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1629394407
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1629394407
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1629394407
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1629394407
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1629394407
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp 1629394407
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1629394407
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_105
timestamp 1629394407
transform 1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1629394407
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1629394407
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1629394407
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1629394407
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1629394407
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1629394407
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1629394407
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1629394407
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1629394407
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1629394407
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1629394407
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1629394407
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1629394407
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp 1629394407
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1629394407
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1629394407
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1629394407
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1629394407
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1629394407
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1629394407
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1629394407
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1629394407
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1629394407
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1629394407
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1629394407
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1629394407
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1629394407
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1629394407
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1629394407
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1629394407
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1629394407
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1629394407
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1629394407
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1629394407
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1629394407
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1629394407
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1629394407
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1629394407
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1629394407
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_105
timestamp 1629394407
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp 1629394407
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1629394407
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1629394407
transform -1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1629394407
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1629394407
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1629394407
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1629394407
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1629394407
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1629394407
transform 1 0 4416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1629394407
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _35_
timestamp 1629394407
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_43
timestamp 1629394407
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1629394407
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1629394407
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 5888 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1629394407
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1629394407
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _31_
timestamp 1629394407
transform 1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_100
timestamp 1629394407
transform 1 0 10304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_88
timestamp 1629394407
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1629394407
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1629394407
transform -1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1629394407
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1629394407
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1629394407
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1629394407
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 4784 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1629394407
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1629394407
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_60
timestamp 1629394407
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1629394407
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _29_
timestamp 1629394407
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1629394407
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _26_
timestamp 1629394407
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1629394407
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1629394407
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp 1629394407
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1629394407
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1629394407
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1629394407
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1629394407
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 3312 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1629394407
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1629394407
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1629394407
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1629394407
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 3956 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1629394407
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 5888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp 1629394407
transform 1 0 6256 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1629394407
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1629394407
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _42_
timestamp 1629394407
transform 1 0 7452 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1629394407
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1629394407
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1629394407
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1629394407
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1629394407
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1629394407
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1629394407
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1629394407
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 2392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1629394407
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _45_
timestamp 1629394407
transform 1 0 4232 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1629394407
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1629394407
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1629394407
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1629394407
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _28_
timestamp 1629394407
transform 1 0 5428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _46_
timestamp 1629394407
transform -1 0 8096 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_76
timestamp 1629394407
transform 1 0 8096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_100
timestamp 1629394407
transform 1 0 10304 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_88
timestamp 1629394407
transform 1 0 9200 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1629394407
transform -1 0 11316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1629394407
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1629394407
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1629394407
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1629394407
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1629394407
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1629394407
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1629394407
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _37_
timestamp 1629394407
transform -1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 4968 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_42
timestamp 1629394407
transform 1 0 4968 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _47_
timestamp 1629394407
transform -1 0 6992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1629394407
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1629394407
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1629394407
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _25_
timestamp 1629394407
transform 1 0 7360 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1629394407
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1629394407
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1629394407
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_105
timestamp 1629394407
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1629394407
transform -1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_11
timestamp 1629394407
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_17
timestamp 1629394407
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1629394407
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1629394407
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1629394407
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1629394407
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1629394407
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _49_
timestamp 1629394407
transform 1 0 2760 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1629394407
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1629394407
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1629394407
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_34
timestamp 1629394407
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1629394407
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform 1 0 4600 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_1  _41_
timestamp 1629394407
transform -1 0 4232 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1629394407
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1629394407
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1629394407
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_46
timestamp 1629394407
transform 1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_54
timestamp 1629394407
transform 1 0 6072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1629394407
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1629394407
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  _24_
timestamp 1629394407
transform 1 0 6348 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1629394407
transform -1 0 8556 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1629394407
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1629394407
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1629394407
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1629394407
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1629394407
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1629394407
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1629394407
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_105
timestamp 1629394407
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1629394407
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1629394407
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1629394407
transform -1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1629394407
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1629394407
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1629394407
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1629394407
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1629394407
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1629394407
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1629394407
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1629394407
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1629394407
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1629394407
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1629394407
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1629394407
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_105
timestamp 1629394407
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1629394407
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1629394407
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1629394407
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1629394407
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1629394407
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1629394407
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1629394407
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1629394407
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1629394407
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1629394407
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1629394407
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1629394407
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1629394407
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1629394407
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1629394407
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_105
timestamp 1629394407
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1629394407
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1629394407
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1629394407
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1629394407
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1629394407
transform -1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp 1629394407
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1629394407
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1629394407
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1629394407
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1629394407
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1629394407
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1629394407
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1629394407
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1629394407
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_81
timestamp 1629394407
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_104
timestamp 1629394407
transform 1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1629394407
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_92
timestamp 1629394407
transform 1 0 9568 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1629394407
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1629394407
transform -1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1629394407
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 5232 11316 5552 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 3600 11316 3920 6 VPWR
port 1 nsew power input
rlabel metal3 s 11635 9800 12435 9920 6 clk
port 2 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 out[0]
port 3 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 out[1]
port 4 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 out[2]
port 5 nsew signal tristate
rlabel metal2 s 2778 13779 2834 14579 6 out[3]
port 6 nsew signal tristate
rlabel metal2 s 9218 13779 9274 14579 6 reset
port 7 nsew signal input
rlabel metal3 s 11635 280 12435 400 6 updown
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12435 14579
<< end >>
